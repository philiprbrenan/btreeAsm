//-----------------------------------------------------------------------------
// Database on a chip synthesis
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree(                                                                      // Test bench for database on a chip
  input                 clock,                                                  // Clock
  input                 reset,                                                  // Reset chip

  input wire [64-1:0] k,
  input wire [8-1:0] d,
  output wire            stop                                            // Program has stopped when this goes high
  );
  integer step;
  integer returnCode;
  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_0_stop||stuckKeys_1_stop||stuckKeys_2_stop||stuckKeys_3_stop||stuckData_0_stop||stuckData_1_stop||stuckData_2_stop||stuckData_3_stop||verilogPut_stop;
  always @ (posedge clock) begin
    if (reset) begin
      step <= -2;
    end
    else begin
      step <= step + 1;
    end
  end
  // process_stuckIsLeaf_0000
  // process_stuckIsFree_0001
  // process_freeNext_0002
  // process_stuckSize_0003
  // process_stuckKeys_0_0004
  // process_stuckKeys_1_0005
  // process_stuckKeys_2_0006
  // process_stuckKeys_3_0007
  // process_stuckData_0_0008
  // process_stuckData_1_0009
  // process_stuckData_2_0010
  // process_stuckData_3_0011
  // process_verilogPut_0012
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[8];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_19_result_0;
  integer stuckIsLeaf_19_requestedAt;
  integer stuckIsLeaf_19_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_19_returnCode;
  integer stuckIsLeaf_20_requestedAt;
  integer stuckIsLeaf_20_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_20_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_19_result_0 <= 0;
      stuckIsLeaf_19_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_19_returnCode <= 0;
      stuckIsLeaf_20_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_20_returnCode <= 0;
      stuckIsLeaf_memory[0] <= 1;
      stuckIsLeaf_memory[1] <= 0;
      stuckIsLeaf_memory[2] <= 0;
      stuckIsLeaf_memory[3] <= 0;
      stuckIsLeaf_memory[4] <= 0;
      stuckIsLeaf_memory[5] <= 0;
      stuckIsLeaf_memory[6] <= 0;
      stuckIsLeaf_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_19_requestedAt > stuckIsLeaf_19_finishedAt && stuckIsLeaf_19_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_19_result_0 <= stuckIsLeaf_memory[verilogPut_stuckIsLeaf_19_index_49];
            stuckIsLeaf_19_finishedAt <= step;
          end
          else if ((stuckIsLeaf_20_requestedAt > stuckIsLeaf_20_finishedAt && stuckIsLeaf_20_requestedAt != step)) begin
            stuckIsLeaf_memory[verilogPut_stuckIsLeaf_20_index_50] <= verilogPut_stuckIsLeaf_20_value_51;
            stuckIsLeaf_20_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[8];
  integer stuckIsFree_23_requestedAt;
  integer stuckIsFree_23_finishedAt;
  integer stuckIsFree_stuckIsFree_23_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_23_finishedAt <= -1;
      stuckIsFree_stuckIsFree_23_returnCode <= 0;
      stuckIsFree_memory[0] <= 0;
      stuckIsFree_memory[1] <= 1;
      stuckIsFree_memory[2] <= 1;
      stuckIsFree_memory[3] <= 1;
      stuckIsFree_memory[4] <= 1;
      stuckIsFree_memory[5] <= 1;
      stuckIsFree_memory[6] <= 1;
      stuckIsFree_memory[7] <= 1;
    end
    else begin                                   // Run the process in full parallel
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_23_requestedAt > stuckIsFree_23_finishedAt && stuckIsFree_23_requestedAt != step)) begin
            stuckIsFree_memory[verilogPut_stuckIsFree_23_index_207] <= verilogPut_stuckIsFree_23_value_208;
            stuckIsFree_23_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [4-1:0] freeNext_memory[8];
  reg [4-1:0] freeNext_freeNext_21_result_0;
  integer freeNext_21_requestedAt;
  integer freeNext_21_finishedAt;
  integer freeNext_freeNext_21_returnCode;
  integer freeNext_22_requestedAt;
  integer freeNext_22_finishedAt;
  integer freeNext_freeNext_22_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_21_result_0 <= 0;
      freeNext_21_finishedAt <= -1;
      freeNext_freeNext_21_returnCode <= 0;
      freeNext_22_finishedAt <= -1;
      freeNext_freeNext_22_returnCode <= 0;
      freeNext_memory[0] <= 1;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 7;
      freeNext_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(freeNext_pc)
        0: begin
          if ((freeNext_21_requestedAt > freeNext_21_finishedAt && freeNext_21_requestedAt != step)) begin
            freeNext_freeNext_21_result_0 <= freeNext_memory[verilogPut_freeNext_21_index_204];
            freeNext_21_finishedAt <= step;
          end
          else if ((freeNext_22_requestedAt > freeNext_22_finishedAt && freeNext_22_requestedAt != step)) begin
            freeNext_memory[verilogPut_freeNext_22_index_205] <= verilogPut_freeNext_22_value_206;
            freeNext_22_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[8];
  reg [3-1:0] stuckSize_stuckSize_17_result_0;
  integer stuckSize_17_requestedAt;
  integer stuckSize_17_finishedAt;
  integer stuckSize_stuckSize_17_returnCode;
  integer stuckSize_18_requestedAt;
  integer stuckSize_18_finishedAt;
  integer stuckSize_stuckSize_18_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_17_result_0 <= 0;
      stuckSize_17_finishedAt <= -1;
      stuckSize_stuckSize_17_returnCode <= 0;
      stuckSize_18_finishedAt <= -1;
      stuckSize_stuckSize_18_returnCode <= 0;
      stuckSize_memory[0] <= 0;
      stuckSize_memory[1] <= 0;
      stuckSize_memory[2] <= 0;
      stuckSize_memory[3] <= 0;
      stuckSize_memory[4] <= 0;
      stuckSize_memory[5] <= 0;
      stuckSize_memory[6] <= 0;
      stuckSize_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_17_requestedAt > stuckSize_17_finishedAt && stuckSize_17_requestedAt != step)) begin
            stuckSize_stuckSize_17_result_0 <= stuckSize_memory[verilogPut_stuckSize_17_index_46];
            stuckSize_17_finishedAt <= step;
          end
          else if ((stuckSize_18_requestedAt > stuckSize_18_finishedAt && stuckSize_18_requestedAt != step)) begin
            stuckSize_memory[verilogPut_stuckSize_18_index_47] <= verilogPut_stuckSize_18_value_48;
            stuckSize_18_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys_0  process_stuckKeys_0_0004
  (* ram_style = "block" *)
  reg [64-1:0] stuckKeys_0_memory[8];
  reg [64-1:0] stuckKeys_0_stuckKeys_0_1_result_0;
  integer stuckKeys_0_1_requestedAt;
  integer stuckKeys_0_1_finishedAt;
  integer stuckKeys_0_stuckKeys_0_1_returnCode;
  integer stuckKeys_0_2_requestedAt;
  integer stuckKeys_0_2_finishedAt;
  integer stuckKeys_0_stuckKeys_0_2_returnCode;
  integer stuckKeys_0_pc;
  integer stuckKeys_0_stop;
  integer stuckKeys_0_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_0_pc <= 0;
      stuckKeys_0_stop <= 0;
      stuckKeys_0_returnCode <= 0;
      stuckKeys_0_stuckKeys_0_1_result_0 <= 0;
      stuckKeys_0_1_finishedAt <= -1;
      stuckKeys_0_stuckKeys_0_1_returnCode <= 0;
      stuckKeys_0_2_finishedAt <= -1;
      stuckKeys_0_stuckKeys_0_2_returnCode <= 0;
      stuckKeys_0_memory[0] <= 0;
      stuckKeys_0_memory[1] <= 0;
      stuckKeys_0_memory[2] <= 0;
      stuckKeys_0_memory[3] <= 0;
      stuckKeys_0_memory[4] <= 0;
      stuckKeys_0_memory[5] <= 0;
      stuckKeys_0_memory[6] <= 0;
      stuckKeys_0_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckKeys_0_pc)
        0: begin
          if ((stuckKeys_0_1_requestedAt > stuckKeys_0_1_finishedAt && stuckKeys_0_1_requestedAt != step)) begin
            stuckKeys_0_stuckKeys_0_1_result_0 <= stuckKeys_0_memory[verilogPut_stuckKeys_0_1_index_10];
            stuckKeys_0_1_finishedAt <= step;
          end
          else if ((stuckKeys_0_2_requestedAt > stuckKeys_0_2_finishedAt && stuckKeys_0_2_requestedAt != step)) begin
            stuckKeys_0_memory[verilogPut_stuckKeys_0_2_index_11] <= verilogPut_stuckKeys_0_2_value_12;
            stuckKeys_0_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_0_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys_1  process_stuckKeys_1_0005
  (* ram_style = "block" *)
  reg [64-1:0] stuckKeys_1_memory[8];
  reg [64-1:0] stuckKeys_1_stuckKeys_1_5_result_0;
  integer stuckKeys_1_5_requestedAt;
  integer stuckKeys_1_5_finishedAt;
  integer stuckKeys_1_stuckKeys_1_5_returnCode;
  integer stuckKeys_1_6_requestedAt;
  integer stuckKeys_1_6_finishedAt;
  integer stuckKeys_1_stuckKeys_1_6_returnCode;
  integer stuckKeys_1_pc;
  integer stuckKeys_1_stop;
  integer stuckKeys_1_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_1_pc <= 0;
      stuckKeys_1_stop <= 0;
      stuckKeys_1_returnCode <= 0;
      stuckKeys_1_stuckKeys_1_5_result_0 <= 0;
      stuckKeys_1_5_finishedAt <= -1;
      stuckKeys_1_stuckKeys_1_5_returnCode <= 0;
      stuckKeys_1_6_finishedAt <= -1;
      stuckKeys_1_stuckKeys_1_6_returnCode <= 0;
      stuckKeys_1_memory[0] <= 0;
      stuckKeys_1_memory[1] <= 0;
      stuckKeys_1_memory[2] <= 0;
      stuckKeys_1_memory[3] <= 0;
      stuckKeys_1_memory[4] <= 0;
      stuckKeys_1_memory[5] <= 0;
      stuckKeys_1_memory[6] <= 0;
      stuckKeys_1_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckKeys_1_pc)
        0: begin
          if ((stuckKeys_1_5_requestedAt > stuckKeys_1_5_finishedAt && stuckKeys_1_5_requestedAt != step)) begin
            stuckKeys_1_stuckKeys_1_5_result_0 <= stuckKeys_1_memory[verilogPut_stuckKeys_1_5_index_20];
            stuckKeys_1_5_finishedAt <= step;
          end
          else if ((stuckKeys_1_6_requestedAt > stuckKeys_1_6_finishedAt && stuckKeys_1_6_requestedAt != step)) begin
            stuckKeys_1_memory[verilogPut_stuckKeys_1_6_index_21] <= verilogPut_stuckKeys_1_6_value_22;
            stuckKeys_1_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_1_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys_2  process_stuckKeys_2_0006
  (* ram_style = "block" *)
  reg [64-1:0] stuckKeys_2_memory[8];
  reg [64-1:0] stuckKeys_2_stuckKeys_2_9_result_0;
  integer stuckKeys_2_9_requestedAt;
  integer stuckKeys_2_9_finishedAt;
  integer stuckKeys_2_stuckKeys_2_9_returnCode;
  integer stuckKeys_2_10_requestedAt;
  integer stuckKeys_2_10_finishedAt;
  integer stuckKeys_2_stuckKeys_2_10_returnCode;
  integer stuckKeys_2_pc;
  integer stuckKeys_2_stop;
  integer stuckKeys_2_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_2_pc <= 0;
      stuckKeys_2_stop <= 0;
      stuckKeys_2_returnCode <= 0;
      stuckKeys_2_stuckKeys_2_9_result_0 <= 0;
      stuckKeys_2_9_finishedAt <= -1;
      stuckKeys_2_stuckKeys_2_9_returnCode <= 0;
      stuckKeys_2_10_finishedAt <= -1;
      stuckKeys_2_stuckKeys_2_10_returnCode <= 0;
      stuckKeys_2_memory[0] <= 0;
      stuckKeys_2_memory[1] <= 0;
      stuckKeys_2_memory[2] <= 0;
      stuckKeys_2_memory[3] <= 0;
      stuckKeys_2_memory[4] <= 0;
      stuckKeys_2_memory[5] <= 0;
      stuckKeys_2_memory[6] <= 0;
      stuckKeys_2_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckKeys_2_pc)
        0: begin
          if ((stuckKeys_2_9_requestedAt > stuckKeys_2_9_finishedAt && stuckKeys_2_9_requestedAt != step)) begin
            stuckKeys_2_stuckKeys_2_9_result_0 <= stuckKeys_2_memory[verilogPut_stuckKeys_2_9_index_30];
            stuckKeys_2_9_finishedAt <= step;
          end
          else if ((stuckKeys_2_10_requestedAt > stuckKeys_2_10_finishedAt && stuckKeys_2_10_requestedAt != step)) begin
            stuckKeys_2_memory[verilogPut_stuckKeys_2_10_index_31] <= verilogPut_stuckKeys_2_10_value_32;
            stuckKeys_2_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_2_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys_3  process_stuckKeys_3_0007
  (* ram_style = "block" *)
  reg [64-1:0] stuckKeys_3_memory[8];
  reg [64-1:0] stuckKeys_3_stuckKeys_3_13_result_0;
  integer stuckKeys_3_13_requestedAt;
  integer stuckKeys_3_13_finishedAt;
  integer stuckKeys_3_stuckKeys_3_13_returnCode;
  integer stuckKeys_3_14_requestedAt;
  integer stuckKeys_3_14_finishedAt;
  integer stuckKeys_3_stuckKeys_3_14_returnCode;
  integer stuckKeys_3_pc;
  integer stuckKeys_3_stop;
  integer stuckKeys_3_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_3_pc <= 0;
      stuckKeys_3_stop <= 0;
      stuckKeys_3_returnCode <= 0;
      stuckKeys_3_stuckKeys_3_13_result_0 <= 0;
      stuckKeys_3_13_finishedAt <= -1;
      stuckKeys_3_stuckKeys_3_13_returnCode <= 0;
      stuckKeys_3_14_finishedAt <= -1;
      stuckKeys_3_stuckKeys_3_14_returnCode <= 0;
      stuckKeys_3_memory[0] <= 0;
      stuckKeys_3_memory[1] <= 0;
      stuckKeys_3_memory[2] <= 0;
      stuckKeys_3_memory[3] <= 0;
      stuckKeys_3_memory[4] <= 0;
      stuckKeys_3_memory[5] <= 0;
      stuckKeys_3_memory[6] <= 0;
      stuckKeys_3_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckKeys_3_pc)
        0: begin
          if ((stuckKeys_3_13_requestedAt > stuckKeys_3_13_finishedAt && stuckKeys_3_13_requestedAt != step)) begin
            stuckKeys_3_stuckKeys_3_13_result_0 <= stuckKeys_3_memory[verilogPut_stuckKeys_3_13_index_40];
            stuckKeys_3_13_finishedAt <= step;
          end
          else if ((stuckKeys_3_14_requestedAt > stuckKeys_3_14_finishedAt && stuckKeys_3_14_requestedAt != step)) begin
            stuckKeys_3_memory[verilogPut_stuckKeys_3_14_index_41] <= verilogPut_stuckKeys_3_14_value_42;
            stuckKeys_3_14_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_3_stop <= 1;
      endcase
    end
  end
  // Process: stuckData_0  process_stuckData_0_0008
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_0_memory[8];
  reg [8-1:0] stuckData_0_stuckData_0_3_result_0;
  integer stuckData_0_3_requestedAt;
  integer stuckData_0_3_finishedAt;
  integer stuckData_0_stuckData_0_3_returnCode;
  integer stuckData_0_4_requestedAt;
  integer stuckData_0_4_finishedAt;
  integer stuckData_0_stuckData_0_4_returnCode;
  integer stuckData_0_pc;
  integer stuckData_0_stop;
  integer stuckData_0_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_0_pc <= 0;
      stuckData_0_stop <= 0;
      stuckData_0_returnCode <= 0;
      stuckData_0_stuckData_0_3_result_0 <= 0;
      stuckData_0_3_finishedAt <= -1;
      stuckData_0_stuckData_0_3_returnCode <= 0;
      stuckData_0_4_finishedAt <= -1;
      stuckData_0_stuckData_0_4_returnCode <= 0;
      stuckData_0_memory[0] <= 0;
      stuckData_0_memory[1] <= 0;
      stuckData_0_memory[2] <= 0;
      stuckData_0_memory[3] <= 0;
      stuckData_0_memory[4] <= 0;
      stuckData_0_memory[5] <= 0;
      stuckData_0_memory[6] <= 0;
      stuckData_0_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckData_0_pc)
        0: begin
          if ((stuckData_0_3_requestedAt > stuckData_0_3_finishedAt && stuckData_0_3_requestedAt != step)) begin
            stuckData_0_stuckData_0_3_result_0 <= stuckData_0_memory[verilogPut_stuckData_0_3_index_13];
            stuckData_0_3_finishedAt <= step;
          end
          else if ((stuckData_0_4_requestedAt > stuckData_0_4_finishedAt && stuckData_0_4_requestedAt != step)) begin
            stuckData_0_memory[verilogPut_stuckData_0_4_index_14] <= verilogPut_stuckData_0_4_value_15;
            stuckData_0_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_0_stop <= 1;
      endcase
    end
  end
  // Process: stuckData_1  process_stuckData_1_0009
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_1_memory[8];
  reg [8-1:0] stuckData_1_stuckData_1_7_result_0;
  integer stuckData_1_7_requestedAt;
  integer stuckData_1_7_finishedAt;
  integer stuckData_1_stuckData_1_7_returnCode;
  integer stuckData_1_8_requestedAt;
  integer stuckData_1_8_finishedAt;
  integer stuckData_1_stuckData_1_8_returnCode;
  integer stuckData_1_pc;
  integer stuckData_1_stop;
  integer stuckData_1_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_1_pc <= 0;
      stuckData_1_stop <= 0;
      stuckData_1_returnCode <= 0;
      stuckData_1_stuckData_1_7_result_0 <= 0;
      stuckData_1_7_finishedAt <= -1;
      stuckData_1_stuckData_1_7_returnCode <= 0;
      stuckData_1_8_finishedAt <= -1;
      stuckData_1_stuckData_1_8_returnCode <= 0;
      stuckData_1_memory[0] <= 0;
      stuckData_1_memory[1] <= 0;
      stuckData_1_memory[2] <= 0;
      stuckData_1_memory[3] <= 0;
      stuckData_1_memory[4] <= 0;
      stuckData_1_memory[5] <= 0;
      stuckData_1_memory[6] <= 0;
      stuckData_1_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckData_1_pc)
        0: begin
          if ((stuckData_1_7_requestedAt > stuckData_1_7_finishedAt && stuckData_1_7_requestedAt != step)) begin
            stuckData_1_stuckData_1_7_result_0 <= stuckData_1_memory[verilogPut_stuckData_1_7_index_23];
            stuckData_1_7_finishedAt <= step;
          end
          else if ((stuckData_1_8_requestedAt > stuckData_1_8_finishedAt && stuckData_1_8_requestedAt != step)) begin
            stuckData_1_memory[verilogPut_stuckData_1_8_index_24] <= verilogPut_stuckData_1_8_value_25;
            stuckData_1_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_1_stop <= 1;
      endcase
    end
  end
  // Process: stuckData_2  process_stuckData_2_0010
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_2_memory[8];
  reg [8-1:0] stuckData_2_stuckData_2_11_result_0;
  integer stuckData_2_11_requestedAt;
  integer stuckData_2_11_finishedAt;
  integer stuckData_2_stuckData_2_11_returnCode;
  integer stuckData_2_12_requestedAt;
  integer stuckData_2_12_finishedAt;
  integer stuckData_2_stuckData_2_12_returnCode;
  integer stuckData_2_pc;
  integer stuckData_2_stop;
  integer stuckData_2_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_2_pc <= 0;
      stuckData_2_stop <= 0;
      stuckData_2_returnCode <= 0;
      stuckData_2_stuckData_2_11_result_0 <= 0;
      stuckData_2_11_finishedAt <= -1;
      stuckData_2_stuckData_2_11_returnCode <= 0;
      stuckData_2_12_finishedAt <= -1;
      stuckData_2_stuckData_2_12_returnCode <= 0;
      stuckData_2_memory[0] <= 0;
      stuckData_2_memory[1] <= 0;
      stuckData_2_memory[2] <= 0;
      stuckData_2_memory[3] <= 0;
      stuckData_2_memory[4] <= 0;
      stuckData_2_memory[5] <= 0;
      stuckData_2_memory[6] <= 0;
      stuckData_2_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckData_2_pc)
        0: begin
          if ((stuckData_2_11_requestedAt > stuckData_2_11_finishedAt && stuckData_2_11_requestedAt != step)) begin
            stuckData_2_stuckData_2_11_result_0 <= stuckData_2_memory[verilogPut_stuckData_2_11_index_33];
            stuckData_2_11_finishedAt <= step;
          end
          else if ((stuckData_2_12_requestedAt > stuckData_2_12_finishedAt && stuckData_2_12_requestedAt != step)) begin
            stuckData_2_memory[verilogPut_stuckData_2_12_index_34] <= verilogPut_stuckData_2_12_value_35;
            stuckData_2_12_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_2_stop <= 1;
      endcase
    end
  end
  // Process: stuckData_3  process_stuckData_3_0011
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_3_memory[8];
  reg [8-1:0] stuckData_3_stuckData_3_15_result_0;
  integer stuckData_3_15_requestedAt;
  integer stuckData_3_15_finishedAt;
  integer stuckData_3_stuckData_3_15_returnCode;
  integer stuckData_3_16_requestedAt;
  integer stuckData_3_16_finishedAt;
  integer stuckData_3_stuckData_3_16_returnCode;
  integer stuckData_3_pc;
  integer stuckData_3_stop;
  integer stuckData_3_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_3_pc <= 0;
      stuckData_3_stop <= 0;
      stuckData_3_returnCode <= 0;
      stuckData_3_stuckData_3_15_result_0 <= 0;
      stuckData_3_15_finishedAt <= -1;
      stuckData_3_stuckData_3_15_returnCode <= 0;
      stuckData_3_16_finishedAt <= -1;
      stuckData_3_stuckData_3_16_returnCode <= 0;
      stuckData_3_memory[0] <= 0;
      stuckData_3_memory[1] <= 0;
      stuckData_3_memory[2] <= 0;
      stuckData_3_memory[3] <= 0;
      stuckData_3_memory[4] <= 0;
      stuckData_3_memory[5] <= 0;
      stuckData_3_memory[6] <= 0;
      stuckData_3_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckData_3_pc)
        0: begin
          if ((stuckData_3_15_requestedAt > stuckData_3_15_finishedAt && stuckData_3_15_requestedAt != step)) begin
            stuckData_3_stuckData_3_15_result_0 <= stuckData_3_memory[verilogPut_stuckData_3_15_index_43];
            stuckData_3_15_finishedAt <= step;
          end
          else if ((stuckData_3_16_requestedAt > stuckData_3_16_finishedAt && stuckData_3_16_requestedAt != step)) begin
            stuckData_3_memory[verilogPut_stuckData_3_16_index_44] <= verilogPut_stuckData_3_16_value_45;
            stuckData_3_16_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_3_stop <= 1;
      endcase
    end
  end
  // Process: verilogPut  process_verilogPut_0012
  reg [64-1:0] verilogPut_k_0;
  reg [8-1:0] verilogPut_d_1;
  reg [4-1:0] verilogPut_index_2;
  reg [3-1:0] verilogPut_size_3;
  reg [1-1:0] verilogPut_isLeaf_4;
  reg [4-1:0] verilogPut_nextFree_5;
  reg [64-1:0] verilogPut_Key_0_6;
  reg [1-1:0] verilogPut_KeyCompares_0_7;
  reg [3-1:0] verilogPut_KeyCollapse_0_8;
  reg [8-1:0] verilogPut_Data_0_9;
  reg [3-1:0] verilogPut_stuckKeys_0_1_index_10;
  reg [3-1:0] verilogPut_stuckKeys_0_2_index_11;
  reg [64-1:0] verilogPut_stuckKeys_0_2_value_12;
  reg [3-1:0] verilogPut_stuckData_0_3_index_13;
  reg [3-1:0] verilogPut_stuckData_0_4_index_14;
  reg [8-1:0] verilogPut_stuckData_0_4_value_15;
  reg [64-1:0] verilogPut_Key_1_16;
  reg [1-1:0] verilogPut_KeyCompares_1_17;
  reg [3-1:0] verilogPut_KeyCollapse_1_18;
  reg [8-1:0] verilogPut_Data_1_19;
  reg [3-1:0] verilogPut_stuckKeys_1_5_index_20;
  reg [3-1:0] verilogPut_stuckKeys_1_6_index_21;
  reg [64-1:0] verilogPut_stuckKeys_1_6_value_22;
  reg [3-1:0] verilogPut_stuckData_1_7_index_23;
  reg [3-1:0] verilogPut_stuckData_1_8_index_24;
  reg [8-1:0] verilogPut_stuckData_1_8_value_25;
  reg [64-1:0] verilogPut_Key_2_26;
  reg [1-1:0] verilogPut_KeyCompares_2_27;
  reg [3-1:0] verilogPut_KeyCollapse_2_28;
  reg [8-1:0] verilogPut_Data_2_29;
  reg [3-1:0] verilogPut_stuckKeys_2_9_index_30;
  reg [3-1:0] verilogPut_stuckKeys_2_10_index_31;
  reg [64-1:0] verilogPut_stuckKeys_2_10_value_32;
  reg [3-1:0] verilogPut_stuckData_2_11_index_33;
  reg [3-1:0] verilogPut_stuckData_2_12_index_34;
  reg [8-1:0] verilogPut_stuckData_2_12_value_35;
  reg [64-1:0] verilogPut_Key_3_36;
  reg [1-1:0] verilogPut_KeyCompares_3_37;
  reg [3-1:0] verilogPut_KeyCollapse_3_38;
  reg [8-1:0] verilogPut_Data_3_39;
  reg [3-1:0] verilogPut_stuckKeys_3_13_index_40;
  reg [3-1:0] verilogPut_stuckKeys_3_14_index_41;
  reg [64-1:0] verilogPut_stuckKeys_3_14_value_42;
  reg [3-1:0] verilogPut_stuckData_3_15_index_43;
  reg [3-1:0] verilogPut_stuckData_3_16_index_44;
  reg [8-1:0] verilogPut_stuckData_3_16_value_45;
  reg [3-1:0] verilogPut_stuckSize_17_index_46;
  reg [3-1:0] verilogPut_stuckSize_18_index_47;
  reg [3-1:0] verilogPut_stuckSize_18_value_48;
  reg [3-1:0] verilogPut_stuckIsLeaf_19_index_49;
  reg [3-1:0] verilogPut_stuckIsLeaf_20_index_50;
  reg [1-1:0] verilogPut_stuckIsLeaf_20_value_51;
  reg [1-1:0] verilogPut_Found_52;
  reg [64-1:0] verilogPut_Key_53;
  reg [64-1:0] verilogPut_FoundKey_54;
  reg [8-1:0] verilogPut_Data_55;
  reg [4-1:0] verilogPut_BtreeIndex_56;
  reg [3-1:0] verilogPut_StuckIndex_57;
  reg [1-1:0] verilogPut_MergeSuccess_58;
  reg [4-1:0] verilogPut_index_59;
  reg [3-1:0] verilogPut_size_60;
  reg [1-1:0] verilogPut_isLeaf_61;
  reg [4-1:0] verilogPut_nextFree_62;
  reg [64-1:0] verilogPut_Key_0_63;
  reg [1-1:0] verilogPut_KeyCompares_0_64;
  reg [3-1:0] verilogPut_KeyCollapse_0_65;
  reg [8-1:0] verilogPut_Data_0_66;
  reg [64-1:0] verilogPut_Key_1_67;
  reg [1-1:0] verilogPut_KeyCompares_1_68;
  reg [3-1:0] verilogPut_KeyCollapse_1_69;
  reg [8-1:0] verilogPut_Data_1_70;
  reg [64-1:0] verilogPut_Key_2_71;
  reg [1-1:0] verilogPut_KeyCompares_2_72;
  reg [3-1:0] verilogPut_KeyCollapse_2_73;
  reg [8-1:0] verilogPut_Data_2_74;
  reg [64-1:0] verilogPut_Key_3_75;
  reg [1-1:0] verilogPut_KeyCompares_3_76;
  reg [3-1:0] verilogPut_KeyCollapse_3_77;
  reg [8-1:0] verilogPut_Data_3_78;
  reg [1-1:0] verilogPut_Found_79;
  reg [64-1:0] verilogPut_Key_80;
  reg [64-1:0] verilogPut_FoundKey_81;
  reg [8-1:0] verilogPut_Data_82;
  reg [4-1:0] verilogPut_BtreeIndex_83;
  reg [3-1:0] verilogPut_StuckIndex_84;
  reg [1-1:0] verilogPut_MergeSuccess_85;
  reg [4-1:0] verilogPut_index_86;
  reg [3-1:0] verilogPut_size_87;
  reg [1-1:0] verilogPut_isLeaf_88;
  reg [4-1:0] verilogPut_nextFree_89;
  reg [64-1:0] verilogPut_Key_0_90;
  reg [1-1:0] verilogPut_KeyCompares_0_91;
  reg [3-1:0] verilogPut_KeyCollapse_0_92;
  reg [8-1:0] verilogPut_Data_0_93;
  reg [64-1:0] verilogPut_Key_1_94;
  reg [1-1:0] verilogPut_KeyCompares_1_95;
  reg [3-1:0] verilogPut_KeyCollapse_1_96;
  reg [8-1:0] verilogPut_Data_1_97;
  reg [64-1:0] verilogPut_Key_2_98;
  reg [1-1:0] verilogPut_KeyCompares_2_99;
  reg [3-1:0] verilogPut_KeyCollapse_2_100;
  reg [8-1:0] verilogPut_Data_2_101;
  reg [64-1:0] verilogPut_Key_3_102;
  reg [1-1:0] verilogPut_KeyCompares_3_103;
  reg [3-1:0] verilogPut_KeyCollapse_3_104;
  reg [8-1:0] verilogPut_Data_3_105;
  reg [1-1:0] verilogPut_Found_106;
  reg [64-1:0] verilogPut_Key_107;
  reg [64-1:0] verilogPut_FoundKey_108;
  reg [8-1:0] verilogPut_Data_109;
  reg [4-1:0] verilogPut_BtreeIndex_110;
  reg [3-1:0] verilogPut_StuckIndex_111;
  reg [1-1:0] verilogPut_MergeSuccess_112;
  reg [4-1:0] verilogPut_child_113;
  reg [4-1:0] verilogPut_parent_114;
  reg [3-1:0] verilogPut_childInparent_115;
  reg [1-1:0] verilogPut_found_116;
  reg [1-1:0] verilogPut_full_117;
  reg [3-1:0] verilogPut_i_118;
  reg [1-1:0] verilogPut_notFull_119;
  reg [4-1:0] verilogPut_index_120;
  reg [3-1:0] verilogPut_size_121;
  reg [1-1:0] verilogPut_isLeaf_122;
  reg [4-1:0] verilogPut_nextFree_123;
  reg [64-1:0] verilogPut_Key_0_124;
  reg [1-1:0] verilogPut_KeyCompares_0_125;
  reg [3-1:0] verilogPut_KeyCollapse_0_126;
  reg [8-1:0] verilogPut_Data_0_127;
  reg [64-1:0] verilogPut_Key_1_128;
  reg [1-1:0] verilogPut_KeyCompares_1_129;
  reg [3-1:0] verilogPut_KeyCollapse_1_130;
  reg [8-1:0] verilogPut_Data_1_131;
  reg [64-1:0] verilogPut_Key_2_132;
  reg [1-1:0] verilogPut_KeyCompares_2_133;
  reg [3-1:0] verilogPut_KeyCollapse_2_134;
  reg [8-1:0] verilogPut_Data_2_135;
  reg [64-1:0] verilogPut_Key_3_136;
  reg [1-1:0] verilogPut_KeyCompares_3_137;
  reg [3-1:0] verilogPut_KeyCollapse_3_138;
  reg [8-1:0] verilogPut_Data_3_139;
  reg [1-1:0] verilogPut_Found_140;
  reg [64-1:0] verilogPut_Key_141;
  reg [64-1:0] verilogPut_FoundKey_142;
  reg [8-1:0] verilogPut_Data_143;
  reg [4-1:0] verilogPut_BtreeIndex_144;
  reg [3-1:0] verilogPut_StuckIndex_145;
  reg [1-1:0] verilogPut_MergeSuccess_146;
  reg [4-1:0] verilogPut_index_147;
  reg [3-1:0] verilogPut_size_148;
  reg [1-1:0] verilogPut_isLeaf_149;
  reg [4-1:0] verilogPut_nextFree_150;
  reg [64-1:0] verilogPut_Key_0_151;
  reg [1-1:0] verilogPut_KeyCompares_0_152;
  reg [3-1:0] verilogPut_KeyCollapse_0_153;
  reg [8-1:0] verilogPut_Data_0_154;
  reg [64-1:0] verilogPut_Key_1_155;
  reg [1-1:0] verilogPut_KeyCompares_1_156;
  reg [3-1:0] verilogPut_KeyCollapse_1_157;
  reg [8-1:0] verilogPut_Data_1_158;
  reg [64-1:0] verilogPut_Key_2_159;
  reg [1-1:0] verilogPut_KeyCompares_2_160;
  reg [3-1:0] verilogPut_KeyCollapse_2_161;
  reg [8-1:0] verilogPut_Data_2_162;
  reg [64-1:0] verilogPut_Key_3_163;
  reg [1-1:0] verilogPut_KeyCompares_3_164;
  reg [3-1:0] verilogPut_KeyCollapse_3_165;
  reg [8-1:0] verilogPut_Data_3_166;
  reg [1-1:0] verilogPut_Found_167;
  reg [64-1:0] verilogPut_Key_168;
  reg [64-1:0] verilogPut_FoundKey_169;
  reg [8-1:0] verilogPut_Data_170;
  reg [4-1:0] verilogPut_BtreeIndex_171;
  reg [3-1:0] verilogPut_StuckIndex_172;
  reg [1-1:0] verilogPut_MergeSuccess_173;
  reg [4-1:0] verilogPut_index_174;
  reg [3-1:0] verilogPut_size_175;
  reg [1-1:0] verilogPut_isLeaf_176;
  reg [4-1:0] verilogPut_nextFree_177;
  reg [64-1:0] verilogPut_Key_0_178;
  reg [1-1:0] verilogPut_KeyCompares_0_179;
  reg [3-1:0] verilogPut_KeyCollapse_0_180;
  reg [8-1:0] verilogPut_Data_0_181;
  reg [64-1:0] verilogPut_Key_1_182;
  reg [1-1:0] verilogPut_KeyCompares_1_183;
  reg [3-1:0] verilogPut_KeyCollapse_1_184;
  reg [8-1:0] verilogPut_Data_1_185;
  reg [64-1:0] verilogPut_Key_2_186;
  reg [1-1:0] verilogPut_KeyCompares_2_187;
  reg [3-1:0] verilogPut_KeyCollapse_2_188;
  reg [8-1:0] verilogPut_Data_2_189;
  reg [64-1:0] verilogPut_Key_3_190;
  reg [1-1:0] verilogPut_KeyCompares_3_191;
  reg [3-1:0] verilogPut_KeyCollapse_3_192;
  reg [8-1:0] verilogPut_Data_3_193;
  reg [1-1:0] verilogPut_Found_194;
  reg [64-1:0] verilogPut_Key_195;
  reg [64-1:0] verilogPut_FoundKey_196;
  reg [8-1:0] verilogPut_Data_197;
  reg [4-1:0] verilogPut_BtreeIndex_198;
  reg [3-1:0] verilogPut_StuckIndex_199;
  reg [1-1:0] verilogPut_MergeSuccess_200;
  reg [4-1:0] verilogPut_indexLeft_201;
  reg [4-1:0] verilogPut_indexRight_202;
  reg [64-1:0] verilogPut_midKey_203;
  reg [3-1:0] verilogPut_freeNext_21_index_204;
  reg [3-1:0] verilogPut_freeNext_22_index_205;
  reg [4-1:0] verilogPut_freeNext_22_value_206;
  reg [3-1:0] verilogPut_stuckIsFree_23_index_207;
  reg [1-1:0] verilogPut_stuckIsFree_23_value_208;
  reg [4-1:0] verilogPut_root_209;
  reg [4-1:0] verilogPut_next_210;
  reg [1-1:0] verilogPut_isLeaf_211;
  reg [1-1:0] verilogPut_isFree_212;
  reg [4-1:0] verilogPut_root_213;
  reg [4-1:0] verilogPut_next_214;
  reg [1-1:0] verilogPut_isLeaf_215;
  reg [1-1:0] verilogPut_isFree_216;
  reg [3-1:0] verilogPut_i_217;
  reg [1-1:0] verilogPut_notFull_218;
  reg [4-1:0] verilogPut_index_219;
  reg [3-1:0] verilogPut_size_220;
  reg [1-1:0] verilogPut_isLeaf_221;
  reg [4-1:0] verilogPut_nextFree_222;
  reg [64-1:0] verilogPut_Key_0_223;
  reg [1-1:0] verilogPut_KeyCompares_0_224;
  reg [3-1:0] verilogPut_KeyCollapse_0_225;
  reg [8-1:0] verilogPut_Data_0_226;
  reg [64-1:0] verilogPut_Key_1_227;
  reg [1-1:0] verilogPut_KeyCompares_1_228;
  reg [3-1:0] verilogPut_KeyCollapse_1_229;
  reg [8-1:0] verilogPut_Data_1_230;
  reg [64-1:0] verilogPut_Key_2_231;
  reg [1-1:0] verilogPut_KeyCompares_2_232;
  reg [3-1:0] verilogPut_KeyCollapse_2_233;
  reg [8-1:0] verilogPut_Data_2_234;
  reg [64-1:0] verilogPut_Key_3_235;
  reg [1-1:0] verilogPut_KeyCompares_3_236;
  reg [3-1:0] verilogPut_KeyCollapse_3_237;
  reg [8-1:0] verilogPut_Data_3_238;
  reg [1-1:0] verilogPut_Found_239;
  reg [64-1:0] verilogPut_Key_240;
  reg [64-1:0] verilogPut_FoundKey_241;
  reg [8-1:0] verilogPut_Data_242;
  reg [4-1:0] verilogPut_BtreeIndex_243;
  reg [3-1:0] verilogPut_StuckIndex_244;
  reg [1-1:0] verilogPut_MergeSuccess_245;
  reg [4-1:0] verilogPut_index_246;
  reg [3-1:0] verilogPut_size_247;
  reg [1-1:0] verilogPut_isLeaf_248;
  reg [4-1:0] verilogPut_nextFree_249;
  reg [64-1:0] verilogPut_Key_0_250;
  reg [1-1:0] verilogPut_KeyCompares_0_251;
  reg [3-1:0] verilogPut_KeyCollapse_0_252;
  reg [8-1:0] verilogPut_Data_0_253;
  reg [64-1:0] verilogPut_Key_1_254;
  reg [1-1:0] verilogPut_KeyCompares_1_255;
  reg [3-1:0] verilogPut_KeyCollapse_1_256;
  reg [8-1:0] verilogPut_Data_1_257;
  reg [64-1:0] verilogPut_Key_2_258;
  reg [1-1:0] verilogPut_KeyCompares_2_259;
  reg [3-1:0] verilogPut_KeyCollapse_2_260;
  reg [8-1:0] verilogPut_Data_2_261;
  reg [64-1:0] verilogPut_Key_3_262;
  reg [1-1:0] verilogPut_KeyCompares_3_263;
  reg [3-1:0] verilogPut_KeyCollapse_3_264;
  reg [8-1:0] verilogPut_Data_3_265;
  reg [1-1:0] verilogPut_Found_266;
  reg [64-1:0] verilogPut_Key_267;
  reg [64-1:0] verilogPut_FoundKey_268;
  reg [8-1:0] verilogPut_Data_269;
  reg [4-1:0] verilogPut_BtreeIndex_270;
  reg [3-1:0] verilogPut_StuckIndex_271;
  reg [1-1:0] verilogPut_MergeSuccess_272;
  reg [4-1:0] verilogPut_index_273;
  reg [3-1:0] verilogPut_size_274;
  reg [1-1:0] verilogPut_isLeaf_275;
  reg [4-1:0] verilogPut_nextFree_276;
  reg [64-1:0] verilogPut_Key_0_277;
  reg [1-1:0] verilogPut_KeyCompares_0_278;
  reg [3-1:0] verilogPut_KeyCollapse_0_279;
  reg [8-1:0] verilogPut_Data_0_280;
  reg [64-1:0] verilogPut_Key_1_281;
  reg [1-1:0] verilogPut_KeyCompares_1_282;
  reg [3-1:0] verilogPut_KeyCollapse_1_283;
  reg [8-1:0] verilogPut_Data_1_284;
  reg [64-1:0] verilogPut_Key_2_285;
  reg [1-1:0] verilogPut_KeyCompares_2_286;
  reg [3-1:0] verilogPut_KeyCollapse_2_287;
  reg [8-1:0] verilogPut_Data_2_288;
  reg [64-1:0] verilogPut_Key_3_289;
  reg [1-1:0] verilogPut_KeyCompares_3_290;
  reg [3-1:0] verilogPut_KeyCollapse_3_291;
  reg [8-1:0] verilogPut_Data_3_292;
  reg [1-1:0] verilogPut_Found_293;
  reg [64-1:0] verilogPut_Key_294;
  reg [64-1:0] verilogPut_FoundKey_295;
  reg [8-1:0] verilogPut_Data_296;
  reg [4-1:0] verilogPut_BtreeIndex_297;
  reg [3-1:0] verilogPut_StuckIndex_298;
  reg [1-1:0] verilogPut_MergeSuccess_299;
  reg [4-1:0] verilogPut_indexLeft_300;
  reg [4-1:0] verilogPut_indexRight_301;
  reg [64-1:0] verilogPut_midKey_302;
  reg [4-1:0] verilogPut_root_303;
  reg [4-1:0] verilogPut_next_304;
  reg [1-1:0] verilogPut_isLeaf_305;
  reg [1-1:0] verilogPut_isFree_306;
  reg [4-1:0] verilogPut_root_307;
  reg [4-1:0] verilogPut_next_308;
  reg [1-1:0] verilogPut_isLeaf_309;
  reg [1-1:0] verilogPut_isFree_310;
  reg [4-1:0] verilogPut_index_311;
  reg [3-1:0] verilogPut_size_312;
  reg [1-1:0] verilogPut_isLeaf_313;
  reg [4-1:0] verilogPut_nextFree_314;
  reg [64-1:0] verilogPut_Key_0_315;
  reg [1-1:0] verilogPut_KeyCompares_0_316;
  reg [3-1:0] verilogPut_KeyCollapse_0_317;
  reg [8-1:0] verilogPut_Data_0_318;
  reg [64-1:0] verilogPut_Key_1_319;
  reg [1-1:0] verilogPut_KeyCompares_1_320;
  reg [3-1:0] verilogPut_KeyCollapse_1_321;
  reg [8-1:0] verilogPut_Data_1_322;
  reg [64-1:0] verilogPut_Key_2_323;
  reg [1-1:0] verilogPut_KeyCompares_2_324;
  reg [3-1:0] verilogPut_KeyCollapse_2_325;
  reg [8-1:0] verilogPut_Data_2_326;
  reg [64-1:0] verilogPut_Key_3_327;
  reg [1-1:0] verilogPut_KeyCompares_3_328;
  reg [3-1:0] verilogPut_KeyCollapse_3_329;
  reg [8-1:0] verilogPut_Data_3_330;
  reg [1-1:0] verilogPut_Found_331;
  reg [64-1:0] verilogPut_Key_332;
  reg [64-1:0] verilogPut_FoundKey_333;
  reg [8-1:0] verilogPut_Data_334;
  reg [4-1:0] verilogPut_BtreeIndex_335;
  reg [3-1:0] verilogPut_StuckIndex_336;
  reg [1-1:0] verilogPut_MergeSuccess_337;
  reg [4-1:0] verilogPut_index_338;
  reg [3-1:0] verilogPut_size_339;
  reg [1-1:0] verilogPut_isLeaf_340;
  reg [4-1:0] verilogPut_nextFree_341;
  reg [64-1:0] verilogPut_Key_0_342;
  reg [1-1:0] verilogPut_KeyCompares_0_343;
  reg [3-1:0] verilogPut_KeyCollapse_0_344;
  reg [8-1:0] verilogPut_Data_0_345;
  reg [64-1:0] verilogPut_Key_1_346;
  reg [1-1:0] verilogPut_KeyCompares_1_347;
  reg [3-1:0] verilogPut_KeyCollapse_1_348;
  reg [8-1:0] verilogPut_Data_1_349;
  reg [64-1:0] verilogPut_Key_2_350;
  reg [1-1:0] verilogPut_KeyCompares_2_351;
  reg [3-1:0] verilogPut_KeyCollapse_2_352;
  reg [8-1:0] verilogPut_Data_2_353;
  reg [64-1:0] verilogPut_Key_3_354;
  reg [1-1:0] verilogPut_KeyCompares_3_355;
  reg [3-1:0] verilogPut_KeyCollapse_3_356;
  reg [8-1:0] verilogPut_Data_3_357;
  reg [1-1:0] verilogPut_Found_358;
  reg [64-1:0] verilogPut_Key_359;
  reg [64-1:0] verilogPut_FoundKey_360;
  reg [8-1:0] verilogPut_Data_361;
  reg [4-1:0] verilogPut_BtreeIndex_362;
  reg [3-1:0] verilogPut_StuckIndex_363;
  reg [1-1:0] verilogPut_MergeSuccess_364;
  reg [4-1:0] verilogPut_index_365;
  reg [3-1:0] verilogPut_size_366;
  reg [1-1:0] verilogPut_isLeaf_367;
  reg [4-1:0] verilogPut_nextFree_368;
  reg [64-1:0] verilogPut_Key_0_369;
  reg [1-1:0] verilogPut_KeyCompares_0_370;
  reg [3-1:0] verilogPut_KeyCollapse_0_371;
  reg [8-1:0] verilogPut_Data_0_372;
  reg [64-1:0] verilogPut_Key_1_373;
  reg [1-1:0] verilogPut_KeyCompares_1_374;
  reg [3-1:0] verilogPut_KeyCollapse_1_375;
  reg [8-1:0] verilogPut_Data_1_376;
  reg [64-1:0] verilogPut_Key_2_377;
  reg [1-1:0] verilogPut_KeyCompares_2_378;
  reg [3-1:0] verilogPut_KeyCollapse_2_379;
  reg [8-1:0] verilogPut_Data_2_380;
  reg [64-1:0] verilogPut_Key_3_381;
  reg [1-1:0] verilogPut_KeyCompares_3_382;
  reg [3-1:0] verilogPut_KeyCollapse_3_383;
  reg [8-1:0] verilogPut_Data_3_384;
  reg [1-1:0] verilogPut_Found_385;
  reg [64-1:0] verilogPut_Key_386;
  reg [64-1:0] verilogPut_FoundKey_387;
  reg [8-1:0] verilogPut_Data_388;
  reg [4-1:0] verilogPut_BtreeIndex_389;
  reg [3-1:0] verilogPut_StuckIndex_390;
  reg [1-1:0] verilogPut_MergeSuccess_391;
  reg [4-1:0] verilogPut_index_392;
  reg [3-1:0] verilogPut_size_393;
  reg [1-1:0] verilogPut_isLeaf_394;
  reg [4-1:0] verilogPut_nextFree_395;
  reg [64-1:0] verilogPut_Key_0_396;
  reg [1-1:0] verilogPut_KeyCompares_0_397;
  reg [3-1:0] verilogPut_KeyCollapse_0_398;
  reg [8-1:0] verilogPut_Data_0_399;
  reg [64-1:0] verilogPut_Key_1_400;
  reg [1-1:0] verilogPut_KeyCompares_1_401;
  reg [3-1:0] verilogPut_KeyCollapse_1_402;
  reg [8-1:0] verilogPut_Data_1_403;
  reg [64-1:0] verilogPut_Key_2_404;
  reg [1-1:0] verilogPut_KeyCompares_2_405;
  reg [3-1:0] verilogPut_KeyCollapse_2_406;
  reg [8-1:0] verilogPut_Data_2_407;
  reg [64-1:0] verilogPut_Key_3_408;
  reg [1-1:0] verilogPut_KeyCompares_3_409;
  reg [3-1:0] verilogPut_KeyCollapse_3_410;
  reg [8-1:0] verilogPut_Data_3_411;
  reg [1-1:0] verilogPut_Found_412;
  reg [64-1:0] verilogPut_Key_413;
  reg [64-1:0] verilogPut_FoundKey_414;
  reg [8-1:0] verilogPut_Data_415;
  reg [4-1:0] verilogPut_BtreeIndex_416;
  reg [3-1:0] verilogPut_StuckIndex_417;
  reg [1-1:0] verilogPut_MergeSuccess_418;
  reg [64-1:0] verilogPut_childKey_419;
  reg [4-1:0] verilogPut_childData_420;
  reg [4-1:0] verilogPut_indexLeft_421;
  reg [4-1:0] verilogPut_indexRight_422;
  reg [64-1:0] verilogPut_midKey_423;
  reg [4-1:0] verilogPut_root_424;
  reg [4-1:0] verilogPut_next_425;
  reg [1-1:0] verilogPut_isLeaf_426;
  reg [1-1:0] verilogPut_isFree_427;
  reg [4-1:0] verilogPut_index_428;
  reg [3-1:0] verilogPut_size_429;
  reg [1-1:0] verilogPut_isLeaf_430;
  reg [4-1:0] verilogPut_nextFree_431;
  reg [64-1:0] verilogPut_Key_0_432;
  reg [1-1:0] verilogPut_KeyCompares_0_433;
  reg [3-1:0] verilogPut_KeyCollapse_0_434;
  reg [8-1:0] verilogPut_Data_0_435;
  reg [64-1:0] verilogPut_Key_1_436;
  reg [1-1:0] verilogPut_KeyCompares_1_437;
  reg [3-1:0] verilogPut_KeyCollapse_1_438;
  reg [8-1:0] verilogPut_Data_1_439;
  reg [64-1:0] verilogPut_Key_2_440;
  reg [1-1:0] verilogPut_KeyCompares_2_441;
  reg [3-1:0] verilogPut_KeyCollapse_2_442;
  reg [8-1:0] verilogPut_Data_2_443;
  reg [64-1:0] verilogPut_Key_3_444;
  reg [1-1:0] verilogPut_KeyCompares_3_445;
  reg [3-1:0] verilogPut_KeyCollapse_3_446;
  reg [8-1:0] verilogPut_Data_3_447;
  reg [1-1:0] verilogPut_Found_448;
  reg [64-1:0] verilogPut_Key_449;
  reg [64-1:0] verilogPut_FoundKey_450;
  reg [8-1:0] verilogPut_Data_451;
  reg [4-1:0] verilogPut_BtreeIndex_452;
  reg [3-1:0] verilogPut_StuckIndex_453;
  reg [1-1:0] verilogPut_MergeSuccess_454;
  reg [4-1:0] verilogPut_index_455;
  reg [3-1:0] verilogPut_size_456;
  reg [1-1:0] verilogPut_isLeaf_457;
  reg [4-1:0] verilogPut_nextFree_458;
  reg [64-1:0] verilogPut_Key_0_459;
  reg [1-1:0] verilogPut_KeyCompares_0_460;
  reg [3-1:0] verilogPut_KeyCollapse_0_461;
  reg [8-1:0] verilogPut_Data_0_462;
  reg [64-1:0] verilogPut_Key_1_463;
  reg [1-1:0] verilogPut_KeyCompares_1_464;
  reg [3-1:0] verilogPut_KeyCollapse_1_465;
  reg [8-1:0] verilogPut_Data_1_466;
  reg [64-1:0] verilogPut_Key_2_467;
  reg [1-1:0] verilogPut_KeyCompares_2_468;
  reg [3-1:0] verilogPut_KeyCollapse_2_469;
  reg [8-1:0] verilogPut_Data_2_470;
  reg [64-1:0] verilogPut_Key_3_471;
  reg [1-1:0] verilogPut_KeyCompares_3_472;
  reg [3-1:0] verilogPut_KeyCollapse_3_473;
  reg [8-1:0] verilogPut_Data_3_474;
  reg [1-1:0] verilogPut_Found_475;
  reg [64-1:0] verilogPut_Key_476;
  reg [64-1:0] verilogPut_FoundKey_477;
  reg [8-1:0] verilogPut_Data_478;
  reg [4-1:0] verilogPut_BtreeIndex_479;
  reg [3-1:0] verilogPut_StuckIndex_480;
  reg [1-1:0] verilogPut_MergeSuccess_481;
  reg [4-1:0] verilogPut_index_482;
  reg [3-1:0] verilogPut_size_483;
  reg [1-1:0] verilogPut_isLeaf_484;
  reg [4-1:0] verilogPut_nextFree_485;
  reg [64-1:0] verilogPut_Key_0_486;
  reg [1-1:0] verilogPut_KeyCompares_0_487;
  reg [3-1:0] verilogPut_KeyCollapse_0_488;
  reg [8-1:0] verilogPut_Data_0_489;
  reg [64-1:0] verilogPut_Key_1_490;
  reg [1-1:0] verilogPut_KeyCompares_1_491;
  reg [3-1:0] verilogPut_KeyCollapse_1_492;
  reg [8-1:0] verilogPut_Data_1_493;
  reg [64-1:0] verilogPut_Key_2_494;
  reg [1-1:0] verilogPut_KeyCompares_2_495;
  reg [3-1:0] verilogPut_KeyCollapse_2_496;
  reg [8-1:0] verilogPut_Data_2_497;
  reg [64-1:0] verilogPut_Key_3_498;
  reg [1-1:0] verilogPut_KeyCompares_3_499;
  reg [3-1:0] verilogPut_KeyCollapse_3_500;
  reg [8-1:0] verilogPut_Data_3_501;
  reg [1-1:0] verilogPut_Found_502;
  reg [64-1:0] verilogPut_Key_503;
  reg [64-1:0] verilogPut_FoundKey_504;
  reg [8-1:0] verilogPut_Data_505;
  reg [4-1:0] verilogPut_BtreeIndex_506;
  reg [3-1:0] verilogPut_StuckIndex_507;
  reg [1-1:0] verilogPut_MergeSuccess_508;
  reg [4-1:0] verilogPut_childIndex_509;
  reg [4-1:0] verilogPut_leftIndex_510;
  reg [64-1:0] verilogPut_midKey_511;
  reg [4-1:0] verilogPut_root_512;
  reg [4-1:0] verilogPut_next_513;
  reg [1-1:0] verilogPut_isLeaf_514;
  reg [1-1:0] verilogPut_isFree_515;
  reg [3-1:0] verilogPut_i_516;
  reg [1-1:0] verilogPut_notFull_517;
  reg [4-1:0] verilogPut_index_518;
  reg [3-1:0] verilogPut_size_519;
  reg [1-1:0] verilogPut_isLeaf_520;
  reg [4-1:0] verilogPut_nextFree_521;
  reg [64-1:0] verilogPut_Key_0_522;
  reg [1-1:0] verilogPut_KeyCompares_0_523;
  reg [3-1:0] verilogPut_KeyCollapse_0_524;
  reg [8-1:0] verilogPut_Data_0_525;
  reg [64-1:0] verilogPut_Key_1_526;
  reg [1-1:0] verilogPut_KeyCompares_1_527;
  reg [3-1:0] verilogPut_KeyCollapse_1_528;
  reg [8-1:0] verilogPut_Data_1_529;
  reg [64-1:0] verilogPut_Key_2_530;
  reg [1-1:0] verilogPut_KeyCompares_2_531;
  reg [3-1:0] verilogPut_KeyCollapse_2_532;
  reg [8-1:0] verilogPut_Data_2_533;
  reg [64-1:0] verilogPut_Key_3_534;
  reg [1-1:0] verilogPut_KeyCompares_3_535;
  reg [3-1:0] verilogPut_KeyCollapse_3_536;
  reg [8-1:0] verilogPut_Data_3_537;
  reg [1-1:0] verilogPut_Found_538;
  reg [64-1:0] verilogPut_Key_539;
  reg [64-1:0] verilogPut_FoundKey_540;
  reg [8-1:0] verilogPut_Data_541;
  reg [4-1:0] verilogPut_BtreeIndex_542;
  reg [3-1:0] verilogPut_StuckIndex_543;
  reg [1-1:0] verilogPut_MergeSuccess_544;
  reg [4-1:0] verilogPut_index_545;
  reg [3-1:0] verilogPut_size_546;
  reg [1-1:0] verilogPut_isLeaf_547;
  reg [4-1:0] verilogPut_nextFree_548;
  reg [64-1:0] verilogPut_Key_0_549;
  reg [1-1:0] verilogPut_KeyCompares_0_550;
  reg [3-1:0] verilogPut_KeyCollapse_0_551;
  reg [8-1:0] verilogPut_Data_0_552;
  reg [64-1:0] verilogPut_Key_1_553;
  reg [1-1:0] verilogPut_KeyCompares_1_554;
  reg [3-1:0] verilogPut_KeyCollapse_1_555;
  reg [8-1:0] verilogPut_Data_1_556;
  reg [64-1:0] verilogPut_Key_2_557;
  reg [1-1:0] verilogPut_KeyCompares_2_558;
  reg [3-1:0] verilogPut_KeyCollapse_2_559;
  reg [8-1:0] verilogPut_Data_2_560;
  reg [64-1:0] verilogPut_Key_3_561;
  reg [1-1:0] verilogPut_KeyCompares_3_562;
  reg [3-1:0] verilogPut_KeyCollapse_3_563;
  reg [8-1:0] verilogPut_Data_3_564;
  reg [1-1:0] verilogPut_Found_565;
  reg [64-1:0] verilogPut_Key_566;
  reg [64-1:0] verilogPut_FoundKey_567;
  reg [8-1:0] verilogPut_Data_568;
  reg [4-1:0] verilogPut_BtreeIndex_569;
  reg [3-1:0] verilogPut_StuckIndex_570;
  reg [1-1:0] verilogPut_MergeSuccess_571;
  reg [4-1:0] verilogPut_index_572;
  reg [3-1:0] verilogPut_size_573;
  reg [1-1:0] verilogPut_isLeaf_574;
  reg [4-1:0] verilogPut_nextFree_575;
  reg [64-1:0] verilogPut_Key_0_576;
  reg [1-1:0] verilogPut_KeyCompares_0_577;
  reg [3-1:0] verilogPut_KeyCollapse_0_578;
  reg [8-1:0] verilogPut_Data_0_579;
  reg [64-1:0] verilogPut_Key_1_580;
  reg [1-1:0] verilogPut_KeyCompares_1_581;
  reg [3-1:0] verilogPut_KeyCollapse_1_582;
  reg [8-1:0] verilogPut_Data_1_583;
  reg [64-1:0] verilogPut_Key_2_584;
  reg [1-1:0] verilogPut_KeyCompares_2_585;
  reg [3-1:0] verilogPut_KeyCollapse_2_586;
  reg [8-1:0] verilogPut_Data_2_587;
  reg [64-1:0] verilogPut_Key_3_588;
  reg [1-1:0] verilogPut_KeyCompares_3_589;
  reg [3-1:0] verilogPut_KeyCollapse_3_590;
  reg [8-1:0] verilogPut_Data_3_591;
  reg [1-1:0] verilogPut_Found_592;
  reg [64-1:0] verilogPut_Key_593;
  reg [64-1:0] verilogPut_FoundKey_594;
  reg [8-1:0] verilogPut_Data_595;
  reg [4-1:0] verilogPut_BtreeIndex_596;
  reg [3-1:0] verilogPut_StuckIndex_597;
  reg [1-1:0] verilogPut_MergeSuccess_598;
  reg [4-1:0] verilogPut_index_599;
  reg [3-1:0] verilogPut_size_600;
  reg [1-1:0] verilogPut_isLeaf_601;
  reg [4-1:0] verilogPut_nextFree_602;
  reg [64-1:0] verilogPut_Key_0_603;
  reg [1-1:0] verilogPut_KeyCompares_0_604;
  reg [3-1:0] verilogPut_KeyCollapse_0_605;
  reg [8-1:0] verilogPut_Data_0_606;
  reg [64-1:0] verilogPut_Key_1_607;
  reg [1-1:0] verilogPut_KeyCompares_1_608;
  reg [3-1:0] verilogPut_KeyCollapse_1_609;
  reg [8-1:0] verilogPut_Data_1_610;
  reg [64-1:0] verilogPut_Key_2_611;
  reg [1-1:0] verilogPut_KeyCompares_2_612;
  reg [3-1:0] verilogPut_KeyCollapse_2_613;
  reg [8-1:0] verilogPut_Data_2_614;
  reg [64-1:0] verilogPut_Key_3_615;
  reg [1-1:0] verilogPut_KeyCompares_3_616;
  reg [3-1:0] verilogPut_KeyCollapse_3_617;
  reg [8-1:0] verilogPut_Data_3_618;
  reg [1-1:0] verilogPut_Found_619;
  reg [64-1:0] verilogPut_Key_620;
  reg [64-1:0] verilogPut_FoundKey_621;
  reg [8-1:0] verilogPut_Data_622;
  reg [4-1:0] verilogPut_BtreeIndex_623;
  reg [3-1:0] verilogPut_StuckIndex_624;
  reg [1-1:0] verilogPut_MergeSuccess_625;
  reg [64-1:0] verilogPut_childKey_626;
  reg [4-1:0] verilogPut_childData_627;
  reg [4-1:0] verilogPut_indexLeft_628;
  reg [4-1:0] verilogPut_indexRight_629;
  reg [64-1:0] verilogPut_midKey_630;
  reg [4-1:0] verilogPut_root_631;
  reg [4-1:0] verilogPut_next_632;
  reg [1-1:0] verilogPut_isLeaf_633;
  reg [1-1:0] verilogPut_isFree_634;
  reg [4-1:0] verilogPut_index_635;
  reg [3-1:0] verilogPut_size_636;
  reg [1-1:0] verilogPut_isLeaf_637;
  reg [4-1:0] verilogPut_nextFree_638;
  reg [64-1:0] verilogPut_Key_0_639;
  reg [1-1:0] verilogPut_KeyCompares_0_640;
  reg [3-1:0] verilogPut_KeyCollapse_0_641;
  reg [8-1:0] verilogPut_Data_0_642;
  reg [64-1:0] verilogPut_Key_1_643;
  reg [1-1:0] verilogPut_KeyCompares_1_644;
  reg [3-1:0] verilogPut_KeyCollapse_1_645;
  reg [8-1:0] verilogPut_Data_1_646;
  reg [64-1:0] verilogPut_Key_2_647;
  reg [1-1:0] verilogPut_KeyCompares_2_648;
  reg [3-1:0] verilogPut_KeyCollapse_2_649;
  reg [8-1:0] verilogPut_Data_2_650;
  reg [64-1:0] verilogPut_Key_3_651;
  reg [1-1:0] verilogPut_KeyCompares_3_652;
  reg [3-1:0] verilogPut_KeyCollapse_3_653;
  reg [8-1:0] verilogPut_Data_3_654;
  reg [1-1:0] verilogPut_Found_655;
  reg [64-1:0] verilogPut_Key_656;
  reg [64-1:0] verilogPut_FoundKey_657;
  reg [8-1:0] verilogPut_Data_658;
  reg [4-1:0] verilogPut_BtreeIndex_659;
  reg [3-1:0] verilogPut_StuckIndex_660;
  reg [1-1:0] verilogPut_MergeSuccess_661;
  reg [4-1:0] verilogPut_index_662;
  reg [3-1:0] verilogPut_size_663;
  reg [1-1:0] verilogPut_isLeaf_664;
  reg [4-1:0] verilogPut_nextFree_665;
  reg [64-1:0] verilogPut_Key_0_666;
  reg [1-1:0] verilogPut_KeyCompares_0_667;
  reg [3-1:0] verilogPut_KeyCollapse_0_668;
  reg [8-1:0] verilogPut_Data_0_669;
  reg [64-1:0] verilogPut_Key_1_670;
  reg [1-1:0] verilogPut_KeyCompares_1_671;
  reg [3-1:0] verilogPut_KeyCollapse_1_672;
  reg [8-1:0] verilogPut_Data_1_673;
  reg [64-1:0] verilogPut_Key_2_674;
  reg [1-1:0] verilogPut_KeyCompares_2_675;
  reg [3-1:0] verilogPut_KeyCollapse_2_676;
  reg [8-1:0] verilogPut_Data_2_677;
  reg [64-1:0] verilogPut_Key_3_678;
  reg [1-1:0] verilogPut_KeyCompares_3_679;
  reg [3-1:0] verilogPut_KeyCollapse_3_680;
  reg [8-1:0] verilogPut_Data_3_681;
  reg [1-1:0] verilogPut_Found_682;
  reg [64-1:0] verilogPut_Key_683;
  reg [64-1:0] verilogPut_FoundKey_684;
  reg [8-1:0] verilogPut_Data_685;
  reg [4-1:0] verilogPut_BtreeIndex_686;
  reg [3-1:0] verilogPut_StuckIndex_687;
  reg [1-1:0] verilogPut_MergeSuccess_688;
  reg [4-1:0] verilogPut_index_689;
  reg [3-1:0] verilogPut_size_690;
  reg [1-1:0] verilogPut_isLeaf_691;
  reg [4-1:0] verilogPut_nextFree_692;
  reg [64-1:0] verilogPut_Key_0_693;
  reg [1-1:0] verilogPut_KeyCompares_0_694;
  reg [3-1:0] verilogPut_KeyCollapse_0_695;
  reg [8-1:0] verilogPut_Data_0_696;
  reg [64-1:0] verilogPut_Key_1_697;
  reg [1-1:0] verilogPut_KeyCompares_1_698;
  reg [3-1:0] verilogPut_KeyCollapse_1_699;
  reg [8-1:0] verilogPut_Data_1_700;
  reg [64-1:0] verilogPut_Key_2_701;
  reg [1-1:0] verilogPut_KeyCompares_2_702;
  reg [3-1:0] verilogPut_KeyCollapse_2_703;
  reg [8-1:0] verilogPut_Data_2_704;
  reg [64-1:0] verilogPut_Key_3_705;
  reg [1-1:0] verilogPut_KeyCompares_3_706;
  reg [3-1:0] verilogPut_KeyCollapse_3_707;
  reg [8-1:0] verilogPut_Data_3_708;
  reg [1-1:0] verilogPut_Found_709;
  reg [64-1:0] verilogPut_Key_710;
  reg [64-1:0] verilogPut_FoundKey_711;
  reg [8-1:0] verilogPut_Data_712;
  reg [4-1:0] verilogPut_BtreeIndex_713;
  reg [3-1:0] verilogPut_StuckIndex_714;
  reg [1-1:0] verilogPut_MergeSuccess_715;
  reg [4-1:0] verilogPut_index_716;
  reg [3-1:0] verilogPut_size_717;
  reg [1-1:0] verilogPut_isLeaf_718;
  reg [4-1:0] verilogPut_nextFree_719;
  reg [64-1:0] verilogPut_Key_0_720;
  reg [1-1:0] verilogPut_KeyCompares_0_721;
  reg [3-1:0] verilogPut_KeyCollapse_0_722;
  reg [8-1:0] verilogPut_Data_0_723;
  reg [64-1:0] verilogPut_Key_1_724;
  reg [1-1:0] verilogPut_KeyCompares_1_725;
  reg [3-1:0] verilogPut_KeyCollapse_1_726;
  reg [8-1:0] verilogPut_Data_1_727;
  reg [64-1:0] verilogPut_Key_2_728;
  reg [1-1:0] verilogPut_KeyCompares_2_729;
  reg [3-1:0] verilogPut_KeyCollapse_2_730;
  reg [8-1:0] verilogPut_Data_2_731;
  reg [64-1:0] verilogPut_Key_3_732;
  reg [1-1:0] verilogPut_KeyCompares_3_733;
  reg [3-1:0] verilogPut_KeyCollapse_3_734;
  reg [8-1:0] verilogPut_Data_3_735;
  reg [1-1:0] verilogPut_Found_736;
  reg [64-1:0] verilogPut_Key_737;
  reg [64-1:0] verilogPut_FoundKey_738;
  reg [8-1:0] verilogPut_Data_739;
  reg [4-1:0] verilogPut_BtreeIndex_740;
  reg [3-1:0] verilogPut_StuckIndex_741;
  reg [1-1:0] verilogPut_MergeSuccess_742;
  reg [64-1:0] verilogPut_childKey_743;
  reg [4-1:0] verilogPut_childData_744;
  reg [4-1:0] verilogPut_indexLeft_745;
  reg [4-1:0] verilogPut_indexRight_746;
  reg [64-1:0] verilogPut_midKey_747;
  reg [4-1:0] verilogPut_root_748;
  reg [4-1:0] verilogPut_next_749;
  reg [1-1:0] verilogPut_isLeaf_750;
  reg [1-1:0] verilogPut_isFree_751;
  reg [4-1:0] verilogPut_index_752;
  reg [3-1:0] verilogPut_size_753;
  reg [1-1:0] verilogPut_isLeaf_754;
  reg [4-1:0] verilogPut_nextFree_755;
  reg [64-1:0] verilogPut_Key_0_756;
  reg [1-1:0] verilogPut_KeyCompares_0_757;
  reg [3-1:0] verilogPut_KeyCollapse_0_758;
  reg [8-1:0] verilogPut_Data_0_759;
  reg [64-1:0] verilogPut_Key_1_760;
  reg [1-1:0] verilogPut_KeyCompares_1_761;
  reg [3-1:0] verilogPut_KeyCollapse_1_762;
  reg [8-1:0] verilogPut_Data_1_763;
  reg [64-1:0] verilogPut_Key_2_764;
  reg [1-1:0] verilogPut_KeyCompares_2_765;
  reg [3-1:0] verilogPut_KeyCollapse_2_766;
  reg [8-1:0] verilogPut_Data_2_767;
  reg [64-1:0] verilogPut_Key_3_768;
  reg [1-1:0] verilogPut_KeyCompares_3_769;
  reg [3-1:0] verilogPut_KeyCollapse_3_770;
  reg [8-1:0] verilogPut_Data_3_771;
  reg [1-1:0] verilogPut_Found_772;
  reg [64-1:0] verilogPut_Key_773;
  reg [64-1:0] verilogPut_FoundKey_774;
  reg [8-1:0] verilogPut_Data_775;
  reg [4-1:0] verilogPut_BtreeIndex_776;
  reg [3-1:0] verilogPut_StuckIndex_777;
  reg [1-1:0] verilogPut_MergeSuccess_778;
  reg [4-1:0] verilogPut_position_779;
  reg [3-1:0] verilogPut_index_780;
  reg [1-1:0] verilogPut_within_781;
  reg [1-1:0] verilogPut_isLeaf_782;
  reg [4-1:0] verilogPut_index_783;
  reg [3-1:0] verilogPut_size_784;
  reg [1-1:0] verilogPut_isLeaf_785;
  reg [4-1:0] verilogPut_nextFree_786;
  reg [64-1:0] verilogPut_Key_0_787;
  reg [1-1:0] verilogPut_KeyCompares_0_788;
  reg [3-1:0] verilogPut_KeyCollapse_0_789;
  reg [8-1:0] verilogPut_Data_0_790;
  reg [64-1:0] verilogPut_Key_1_791;
  reg [1-1:0] verilogPut_KeyCompares_1_792;
  reg [3-1:0] verilogPut_KeyCollapse_1_793;
  reg [8-1:0] verilogPut_Data_1_794;
  reg [64-1:0] verilogPut_Key_2_795;
  reg [1-1:0] verilogPut_KeyCompares_2_796;
  reg [3-1:0] verilogPut_KeyCollapse_2_797;
  reg [8-1:0] verilogPut_Data_2_798;
  reg [64-1:0] verilogPut_Key_3_799;
  reg [1-1:0] verilogPut_KeyCompares_3_800;
  reg [3-1:0] verilogPut_KeyCollapse_3_801;
  reg [8-1:0] verilogPut_Data_3_802;
  reg [1-1:0] verilogPut_Found_803;
  reg [64-1:0] verilogPut_Key_804;
  reg [64-1:0] verilogPut_FoundKey_805;
  reg [8-1:0] verilogPut_Data_806;
  reg [4-1:0] verilogPut_BtreeIndex_807;
  reg [3-1:0] verilogPut_StuckIndex_808;
  reg [1-1:0] verilogPut_MergeSuccess_809;
  reg [4-1:0] verilogPut_index_810;
  reg [3-1:0] verilogPut_size_811;
  reg [1-1:0] verilogPut_isLeaf_812;
  reg [4-1:0] verilogPut_nextFree_813;
  reg [64-1:0] verilogPut_Key_0_814;
  reg [1-1:0] verilogPut_KeyCompares_0_815;
  reg [3-1:0] verilogPut_KeyCollapse_0_816;
  reg [8-1:0] verilogPut_Data_0_817;
  reg [64-1:0] verilogPut_Key_1_818;
  reg [1-1:0] verilogPut_KeyCompares_1_819;
  reg [3-1:0] verilogPut_KeyCollapse_1_820;
  reg [8-1:0] verilogPut_Data_1_821;
  reg [64-1:0] verilogPut_Key_2_822;
  reg [1-1:0] verilogPut_KeyCompares_2_823;
  reg [3-1:0] verilogPut_KeyCollapse_2_824;
  reg [8-1:0] verilogPut_Data_2_825;
  reg [64-1:0] verilogPut_Key_3_826;
  reg [1-1:0] verilogPut_KeyCompares_3_827;
  reg [3-1:0] verilogPut_KeyCollapse_3_828;
  reg [8-1:0] verilogPut_Data_3_829;
  reg [1-1:0] verilogPut_Found_830;
  reg [64-1:0] verilogPut_Key_831;
  reg [64-1:0] verilogPut_FoundKey_832;
  reg [8-1:0] verilogPut_Data_833;
  reg [4-1:0] verilogPut_BtreeIndex_834;
  reg [3-1:0] verilogPut_StuckIndex_835;
  reg [1-1:0] verilogPut_MergeSuccess_836;
  reg [4-1:0] verilogPut_index_837;
  reg [3-1:0] verilogPut_size_838;
  reg [1-1:0] verilogPut_isLeaf_839;
  reg [4-1:0] verilogPut_nextFree_840;
  reg [64-1:0] verilogPut_Key_0_841;
  reg [1-1:0] verilogPut_KeyCompares_0_842;
  reg [3-1:0] verilogPut_KeyCollapse_0_843;
  reg [8-1:0] verilogPut_Data_0_844;
  reg [64-1:0] verilogPut_Key_1_845;
  reg [1-1:0] verilogPut_KeyCompares_1_846;
  reg [3-1:0] verilogPut_KeyCollapse_1_847;
  reg [8-1:0] verilogPut_Data_1_848;
  reg [64-1:0] verilogPut_Key_2_849;
  reg [1-1:0] verilogPut_KeyCompares_2_850;
  reg [3-1:0] verilogPut_KeyCollapse_2_851;
  reg [8-1:0] verilogPut_Data_2_852;
  reg [64-1:0] verilogPut_Key_3_853;
  reg [1-1:0] verilogPut_KeyCompares_3_854;
  reg [3-1:0] verilogPut_KeyCollapse_3_855;
  reg [8-1:0] verilogPut_Data_3_856;
  reg [1-1:0] verilogPut_Found_857;
  reg [64-1:0] verilogPut_Key_858;
  reg [64-1:0] verilogPut_FoundKey_859;
  reg [8-1:0] verilogPut_Data_860;
  reg [4-1:0] verilogPut_BtreeIndex_861;
  reg [3-1:0] verilogPut_StuckIndex_862;
  reg [1-1:0] verilogPut_MergeSuccess_863;
  reg [64-1:0] verilogPut_childKey_864;
  reg [4-1:0] verilogPut_childData_865;
  reg [4-1:0] verilogPut_indexLeft_866;
  reg [4-1:0] verilogPut_indexRight_867;
  reg [64-1:0] verilogPut_midKey_868;
  reg [1-1:0] verilogPut_success_869;
  reg [1-1:0] verilogPut_test_870;
  reg [4-1:0] verilogPut_next_871;
  reg [4-1:0] verilogPut_root_872;
  reg [1-1:0] verilogPut_isFree_873;
  reg [4-1:0] verilogPut_next_874;
  reg [4-1:0] verilogPut_root_875;
  reg [1-1:0] verilogPut_isFree_876;
  reg [4-1:0] verilogPut_index_877;
  reg [3-1:0] verilogPut_size_878;
  reg [1-1:0] verilogPut_isLeaf_879;
  reg [4-1:0] verilogPut_nextFree_880;
  reg [64-1:0] verilogPut_Key_0_881;
  reg [1-1:0] verilogPut_KeyCompares_0_882;
  reg [3-1:0] verilogPut_KeyCollapse_0_883;
  reg [8-1:0] verilogPut_Data_0_884;
  reg [64-1:0] verilogPut_Key_1_885;
  reg [1-1:0] verilogPut_KeyCompares_1_886;
  reg [3-1:0] verilogPut_KeyCollapse_1_887;
  reg [8-1:0] verilogPut_Data_1_888;
  reg [64-1:0] verilogPut_Key_2_889;
  reg [1-1:0] verilogPut_KeyCompares_2_890;
  reg [3-1:0] verilogPut_KeyCollapse_2_891;
  reg [8-1:0] verilogPut_Data_2_892;
  reg [64-1:0] verilogPut_Key_3_893;
  reg [1-1:0] verilogPut_KeyCompares_3_894;
  reg [3-1:0] verilogPut_KeyCollapse_3_895;
  reg [8-1:0] verilogPut_Data_3_896;
  reg [1-1:0] verilogPut_Found_897;
  reg [64-1:0] verilogPut_Key_898;
  reg [64-1:0] verilogPut_FoundKey_899;
  reg [8-1:0] verilogPut_Data_900;
  reg [4-1:0] verilogPut_BtreeIndex_901;
  reg [3-1:0] verilogPut_StuckIndex_902;
  reg [1-1:0] verilogPut_MergeSuccess_903;
  reg [4-1:0] verilogPut_index_904;
  reg [3-1:0] verilogPut_size_905;
  reg [1-1:0] verilogPut_isLeaf_906;
  reg [4-1:0] verilogPut_nextFree_907;
  reg [64-1:0] verilogPut_Key_0_908;
  reg [1-1:0] verilogPut_KeyCompares_0_909;
  reg [3-1:0] verilogPut_KeyCollapse_0_910;
  reg [8-1:0] verilogPut_Data_0_911;
  reg [64-1:0] verilogPut_Key_1_912;
  reg [1-1:0] verilogPut_KeyCompares_1_913;
  reg [3-1:0] verilogPut_KeyCollapse_1_914;
  reg [8-1:0] verilogPut_Data_1_915;
  reg [64-1:0] verilogPut_Key_2_916;
  reg [1-1:0] verilogPut_KeyCompares_2_917;
  reg [3-1:0] verilogPut_KeyCollapse_2_918;
  reg [8-1:0] verilogPut_Data_2_919;
  reg [64-1:0] verilogPut_Key_3_920;
  reg [1-1:0] verilogPut_KeyCompares_3_921;
  reg [3-1:0] verilogPut_KeyCollapse_3_922;
  reg [8-1:0] verilogPut_Data_3_923;
  reg [1-1:0] verilogPut_Found_924;
  reg [64-1:0] verilogPut_Key_925;
  reg [64-1:0] verilogPut_FoundKey_926;
  reg [8-1:0] verilogPut_Data_927;
  reg [4-1:0] verilogPut_BtreeIndex_928;
  reg [3-1:0] verilogPut_StuckIndex_929;
  reg [1-1:0] verilogPut_MergeSuccess_930;
  reg [4-1:0] verilogPut_index_931;
  reg [3-1:0] verilogPut_size_932;
  reg [1-1:0] verilogPut_isLeaf_933;
  reg [4-1:0] verilogPut_nextFree_934;
  reg [64-1:0] verilogPut_Key_0_935;
  reg [1-1:0] verilogPut_KeyCompares_0_936;
  reg [3-1:0] verilogPut_KeyCollapse_0_937;
  reg [8-1:0] verilogPut_Data_0_938;
  reg [64-1:0] verilogPut_Key_1_939;
  reg [1-1:0] verilogPut_KeyCompares_1_940;
  reg [3-1:0] verilogPut_KeyCollapse_1_941;
  reg [8-1:0] verilogPut_Data_1_942;
  reg [64-1:0] verilogPut_Key_2_943;
  reg [1-1:0] verilogPut_KeyCompares_2_944;
  reg [3-1:0] verilogPut_KeyCollapse_2_945;
  reg [8-1:0] verilogPut_Data_2_946;
  reg [64-1:0] verilogPut_Key_3_947;
  reg [1-1:0] verilogPut_KeyCompares_3_948;
  reg [3-1:0] verilogPut_KeyCollapse_3_949;
  reg [8-1:0] verilogPut_Data_3_950;
  reg [1-1:0] verilogPut_Found_951;
  reg [64-1:0] verilogPut_Key_952;
  reg [64-1:0] verilogPut_FoundKey_953;
  reg [8-1:0] verilogPut_Data_954;
  reg [4-1:0] verilogPut_BtreeIndex_955;
  reg [3-1:0] verilogPut_StuckIndex_956;
  reg [1-1:0] verilogPut_MergeSuccess_957;
  reg [64-1:0] verilogPut_childKey_958;
  reg [3-1:0] verilogPut_leftChild_959;
  reg [3-1:0] verilogPut_rightChild_960;
  reg [4-1:0] verilogPut_childData_961;
  reg [4-1:0] verilogPut_indexLeft_962;
  reg [4-1:0] verilogPut_indexRight_963;
  reg [64-1:0] verilogPut_midKey_964;
  reg [1-1:0] verilogPut_success_965;
  reg [1-1:0] verilogPut_test_966;
  reg [4-1:0] verilogPut_next_967;
  reg [4-1:0] verilogPut_root_968;
  reg [1-1:0] verilogPut_isFree_969;
  reg [4-1:0] verilogPut_next_970;
  reg [4-1:0] verilogPut_root_971;
  reg [1-1:0] verilogPut_isFree_972;
  reg [4-1:0] verilogPut_index_973;
  reg [3-1:0] verilogPut_size_974;
  reg [1-1:0] verilogPut_isLeaf_975;
  reg [4-1:0] verilogPut_nextFree_976;
  reg [64-1:0] verilogPut_Key_0_977;
  reg [1-1:0] verilogPut_KeyCompares_0_978;
  reg [3-1:0] verilogPut_KeyCollapse_0_979;
  reg [8-1:0] verilogPut_Data_0_980;
  reg [64-1:0] verilogPut_Key_1_981;
  reg [1-1:0] verilogPut_KeyCompares_1_982;
  reg [3-1:0] verilogPut_KeyCollapse_1_983;
  reg [8-1:0] verilogPut_Data_1_984;
  reg [64-1:0] verilogPut_Key_2_985;
  reg [1-1:0] verilogPut_KeyCompares_2_986;
  reg [3-1:0] verilogPut_KeyCollapse_2_987;
  reg [8-1:0] verilogPut_Data_2_988;
  reg [64-1:0] verilogPut_Key_3_989;
  reg [1-1:0] verilogPut_KeyCompares_3_990;
  reg [3-1:0] verilogPut_KeyCollapse_3_991;
  reg [8-1:0] verilogPut_Data_3_992;
  reg [1-1:0] verilogPut_Found_993;
  reg [64-1:0] verilogPut_Key_994;
  reg [64-1:0] verilogPut_FoundKey_995;
  reg [8-1:0] verilogPut_Data_996;
  reg [4-1:0] verilogPut_BtreeIndex_997;
  reg [3-1:0] verilogPut_StuckIndex_998;
  reg [1-1:0] verilogPut_MergeSuccess_999;
  reg [4-1:0] verilogPut_index_1000;
  reg [3-1:0] verilogPut_size_1001;
  reg [1-1:0] verilogPut_isLeaf_1002;
  reg [4-1:0] verilogPut_nextFree_1003;
  reg [64-1:0] verilogPut_Key_0_1004;
  reg [1-1:0] verilogPut_KeyCompares_0_1005;
  reg [3-1:0] verilogPut_KeyCollapse_0_1006;
  reg [8-1:0] verilogPut_Data_0_1007;
  reg [64-1:0] verilogPut_Key_1_1008;
  reg [1-1:0] verilogPut_KeyCompares_1_1009;
  reg [3-1:0] verilogPut_KeyCollapse_1_1010;
  reg [8-1:0] verilogPut_Data_1_1011;
  reg [64-1:0] verilogPut_Key_2_1012;
  reg [1-1:0] verilogPut_KeyCompares_2_1013;
  reg [3-1:0] verilogPut_KeyCollapse_2_1014;
  reg [8-1:0] verilogPut_Data_2_1015;
  reg [64-1:0] verilogPut_Key_3_1016;
  reg [1-1:0] verilogPut_KeyCompares_3_1017;
  reg [3-1:0] verilogPut_KeyCollapse_3_1018;
  reg [8-1:0] verilogPut_Data_3_1019;
  reg [1-1:0] verilogPut_Found_1020;
  reg [64-1:0] verilogPut_Key_1021;
  reg [64-1:0] verilogPut_FoundKey_1022;
  reg [8-1:0] verilogPut_Data_1023;
  reg [4-1:0] verilogPut_BtreeIndex_1024;
  reg [3-1:0] verilogPut_StuckIndex_1025;
  reg [1-1:0] verilogPut_MergeSuccess_1026;
  reg [64-1:0] verilogPut_childKey_1027;
  reg [3-1:0] verilogPut_size_1028;
  reg [4-1:0] verilogPut_childData_1029;
  reg [4-1:0] verilogPut_indexLeft_1030;
  reg [4-1:0] verilogPut_indexRight_1031;
  reg [64-1:0] verilogPut_midKey_1032;
  reg [1-1:0] verilogPut_success_1033;
  reg [1-1:0] verilogPut_test_1034;
  reg [4-1:0] verilogPut_next_1035;
  reg [4-1:0] verilogPut_root_1036;
  reg [1-1:0] verilogPut_isFree_1037;
  reg [4-1:0] verilogPut_index_1038;
  reg [3-1:0] verilogPut_size_1039;
  reg [1-1:0] verilogPut_isLeaf_1040;
  reg [4-1:0] verilogPut_nextFree_1041;
  reg [64-1:0] verilogPut_Key_0_1042;
  reg [1-1:0] verilogPut_KeyCompares_0_1043;
  reg [3-1:0] verilogPut_KeyCollapse_0_1044;
  reg [8-1:0] verilogPut_Data_0_1045;
  reg [64-1:0] verilogPut_Key_1_1046;
  reg [1-1:0] verilogPut_KeyCompares_1_1047;
  reg [3-1:0] verilogPut_KeyCollapse_1_1048;
  reg [8-1:0] verilogPut_Data_1_1049;
  reg [64-1:0] verilogPut_Key_2_1050;
  reg [1-1:0] verilogPut_KeyCompares_2_1051;
  reg [3-1:0] verilogPut_KeyCollapse_2_1052;
  reg [8-1:0] verilogPut_Data_2_1053;
  reg [64-1:0] verilogPut_Key_3_1054;
  reg [1-1:0] verilogPut_KeyCompares_3_1055;
  reg [3-1:0] verilogPut_KeyCollapse_3_1056;
  reg [8-1:0] verilogPut_Data_3_1057;
  reg [1-1:0] verilogPut_Found_1058;
  reg [64-1:0] verilogPut_Key_1059;
  reg [64-1:0] verilogPut_FoundKey_1060;
  reg [8-1:0] verilogPut_Data_1061;
  reg [4-1:0] verilogPut_BtreeIndex_1062;
  reg [3-1:0] verilogPut_StuckIndex_1063;
  reg [1-1:0] verilogPut_MergeSuccess_1064;
  reg [4-1:0] verilogPut_index_1065;
  reg [3-1:0] verilogPut_size_1066;
  reg [1-1:0] verilogPut_isLeaf_1067;
  reg [4-1:0] verilogPut_nextFree_1068;
  reg [64-1:0] verilogPut_Key_0_1069;
  reg [1-1:0] verilogPut_KeyCompares_0_1070;
  reg [3-1:0] verilogPut_KeyCollapse_0_1071;
  reg [8-1:0] verilogPut_Data_0_1072;
  reg [64-1:0] verilogPut_Key_1_1073;
  reg [1-1:0] verilogPut_KeyCompares_1_1074;
  reg [3-1:0] verilogPut_KeyCollapse_1_1075;
  reg [8-1:0] verilogPut_Data_1_1076;
  reg [64-1:0] verilogPut_Key_2_1077;
  reg [1-1:0] verilogPut_KeyCompares_2_1078;
  reg [3-1:0] verilogPut_KeyCollapse_2_1079;
  reg [8-1:0] verilogPut_Data_2_1080;
  reg [64-1:0] verilogPut_Key_3_1081;
  reg [1-1:0] verilogPut_KeyCompares_3_1082;
  reg [3-1:0] verilogPut_KeyCollapse_3_1083;
  reg [8-1:0] verilogPut_Data_3_1084;
  reg [1-1:0] verilogPut_Found_1085;
  reg [64-1:0] verilogPut_Key_1086;
  reg [64-1:0] verilogPut_FoundKey_1087;
  reg [8-1:0] verilogPut_Data_1088;
  reg [4-1:0] verilogPut_BtreeIndex_1089;
  reg [3-1:0] verilogPut_StuckIndex_1090;
  reg [1-1:0] verilogPut_MergeSuccess_1091;
  reg [64-1:0] verilogPut_childKey_1092;
  reg [3-1:0] verilogPut_size_1093;
  reg [4-1:0] verilogPut_childData_1094;
  reg [4-1:0] verilogPut_indexLeft_1095;
  reg [4-1:0] verilogPut_indexRight_1096;
  reg [64-1:0] verilogPut_midKey_1097;
  reg [1-1:0] verilogPut_success_1098;
  reg [1-1:0] verilogPut_test_1099;
  reg [4-1:0] verilogPut_next_1100;
  reg [4-1:0] verilogPut_root_1101;
  reg [1-1:0] verilogPut_isFree_1102;
  reg [4-1:0] verilogPut_index_1103;
  reg [3-1:0] verilogPut_size_1104;
  reg [1-1:0] verilogPut_isLeaf_1105;
  reg [4-1:0] verilogPut_nextFree_1106;
  reg [64-1:0] verilogPut_Key_0_1107;
  reg [1-1:0] verilogPut_KeyCompares_0_1108;
  reg [3-1:0] verilogPut_KeyCollapse_0_1109;
  reg [8-1:0] verilogPut_Data_0_1110;
  reg [64-1:0] verilogPut_Key_1_1111;
  reg [1-1:0] verilogPut_KeyCompares_1_1112;
  reg [3-1:0] verilogPut_KeyCollapse_1_1113;
  reg [8-1:0] verilogPut_Data_1_1114;
  reg [64-1:0] verilogPut_Key_2_1115;
  reg [1-1:0] verilogPut_KeyCompares_2_1116;
  reg [3-1:0] verilogPut_KeyCollapse_2_1117;
  reg [8-1:0] verilogPut_Data_2_1118;
  reg [64-1:0] verilogPut_Key_3_1119;
  reg [1-1:0] verilogPut_KeyCompares_3_1120;
  reg [3-1:0] verilogPut_KeyCollapse_3_1121;
  reg [8-1:0] verilogPut_Data_3_1122;
  reg [1-1:0] verilogPut_Found_1123;
  reg [64-1:0] verilogPut_Key_1124;
  reg [64-1:0] verilogPut_FoundKey_1125;
  reg [8-1:0] verilogPut_Data_1126;
  reg [4-1:0] verilogPut_BtreeIndex_1127;
  reg [3-1:0] verilogPut_StuckIndex_1128;
  reg [1-1:0] verilogPut_MergeSuccess_1129;
  reg [4-1:0] verilogPut_index_1130;
  reg [3-1:0] verilogPut_size_1131;
  reg [1-1:0] verilogPut_isLeaf_1132;
  reg [4-1:0] verilogPut_nextFree_1133;
  reg [64-1:0] verilogPut_Key_0_1134;
  reg [1-1:0] verilogPut_KeyCompares_0_1135;
  reg [3-1:0] verilogPut_KeyCollapse_0_1136;
  reg [8-1:0] verilogPut_Data_0_1137;
  reg [64-1:0] verilogPut_Key_1_1138;
  reg [1-1:0] verilogPut_KeyCompares_1_1139;
  reg [3-1:0] verilogPut_KeyCollapse_1_1140;
  reg [8-1:0] verilogPut_Data_1_1141;
  reg [64-1:0] verilogPut_Key_2_1142;
  reg [1-1:0] verilogPut_KeyCompares_2_1143;
  reg [3-1:0] verilogPut_KeyCollapse_2_1144;
  reg [8-1:0] verilogPut_Data_2_1145;
  reg [64-1:0] verilogPut_Key_3_1146;
  reg [1-1:0] verilogPut_KeyCompares_3_1147;
  reg [3-1:0] verilogPut_KeyCollapse_3_1148;
  reg [8-1:0] verilogPut_Data_3_1149;
  reg [1-1:0] verilogPut_Found_1150;
  reg [64-1:0] verilogPut_Key_1151;
  reg [64-1:0] verilogPut_FoundKey_1152;
  reg [8-1:0] verilogPut_Data_1153;
  reg [4-1:0] verilogPut_BtreeIndex_1154;
  reg [3-1:0] verilogPut_StuckIndex_1155;
  reg [1-1:0] verilogPut_MergeSuccess_1156;
  reg [64-1:0] verilogPut_childKey_1157;
  reg [4-1:0] verilogPut_childData_1158;
  reg [4-1:0] verilogPut_indexLeft_1159;
  reg [4-1:0] verilogPut_indexRight_1160;
  reg [64-1:0] verilogPut_midKey_1161;
  reg [1-1:0] verilogPut_success_1162;
  reg [1-1:0] verilogPut_test_1163;
  reg [4-1:0] verilogPut_next_1164;
  reg [4-1:0] verilogPut_root_1165;
  reg [1-1:0] verilogPut_isFree_1166;
  reg [4-1:0] verilogPut_index_1167;
  reg [3-1:0] verilogPut_size_1168;
  reg [1-1:0] verilogPut_isLeaf_1169;
  reg [4-1:0] verilogPut_nextFree_1170;
  reg [64-1:0] verilogPut_Key_0_1171;
  reg [1-1:0] verilogPut_KeyCompares_0_1172;
  reg [3-1:0] verilogPut_KeyCollapse_0_1173;
  reg [8-1:0] verilogPut_Data_0_1174;
  reg [64-1:0] verilogPut_Key_1_1175;
  reg [1-1:0] verilogPut_KeyCompares_1_1176;
  reg [3-1:0] verilogPut_KeyCollapse_1_1177;
  reg [8-1:0] verilogPut_Data_1_1178;
  reg [64-1:0] verilogPut_Key_2_1179;
  reg [1-1:0] verilogPut_KeyCompares_2_1180;
  reg [3-1:0] verilogPut_KeyCollapse_2_1181;
  reg [8-1:0] verilogPut_Data_2_1182;
  reg [64-1:0] verilogPut_Key_3_1183;
  reg [1-1:0] verilogPut_KeyCompares_3_1184;
  reg [3-1:0] verilogPut_KeyCollapse_3_1185;
  reg [8-1:0] verilogPut_Data_3_1186;
  reg [1-1:0] verilogPut_Found_1187;
  reg [64-1:0] verilogPut_Key_1188;
  reg [64-1:0] verilogPut_FoundKey_1189;
  reg [8-1:0] verilogPut_Data_1190;
  reg [4-1:0] verilogPut_BtreeIndex_1191;
  reg [3-1:0] verilogPut_StuckIndex_1192;
  reg [1-1:0] verilogPut_MergeSuccess_1193;
  reg [4-1:0] verilogPut_index_1194;
  reg [3-1:0] verilogPut_size_1195;
  reg [1-1:0] verilogPut_isLeaf_1196;
  reg [4-1:0] verilogPut_nextFree_1197;
  reg [64-1:0] verilogPut_Key_0_1198;
  reg [1-1:0] verilogPut_KeyCompares_0_1199;
  reg [3-1:0] verilogPut_KeyCollapse_0_1200;
  reg [8-1:0] verilogPut_Data_0_1201;
  reg [64-1:0] verilogPut_Key_1_1202;
  reg [1-1:0] verilogPut_KeyCompares_1_1203;
  reg [3-1:0] verilogPut_KeyCollapse_1_1204;
  reg [8-1:0] verilogPut_Data_1_1205;
  reg [64-1:0] verilogPut_Key_2_1206;
  reg [1-1:0] verilogPut_KeyCompares_2_1207;
  reg [3-1:0] verilogPut_KeyCollapse_2_1208;
  reg [8-1:0] verilogPut_Data_2_1209;
  reg [64-1:0] verilogPut_Key_3_1210;
  reg [1-1:0] verilogPut_KeyCompares_3_1211;
  reg [3-1:0] verilogPut_KeyCollapse_3_1212;
  reg [8-1:0] verilogPut_Data_3_1213;
  reg [1-1:0] verilogPut_Found_1214;
  reg [64-1:0] verilogPut_Key_1215;
  reg [64-1:0] verilogPut_FoundKey_1216;
  reg [8-1:0] verilogPut_Data_1217;
  reg [4-1:0] verilogPut_BtreeIndex_1218;
  reg [3-1:0] verilogPut_StuckIndex_1219;
  reg [1-1:0] verilogPut_MergeSuccess_1220;
  reg [64-1:0] verilogPut_childKey_1221;
  reg [3-1:0] verilogPut_leftChild_1222;
  reg [3-1:0] verilogPut_rightChild_1223;
  reg [4-1:0] verilogPut_childData_1224;
  reg [4-1:0] verilogPut_indexLeft_1225;
  reg [4-1:0] verilogPut_indexRight_1226;
  reg [64-1:0] verilogPut_midKey_1227;
  reg [1-1:0] verilogPut_success_1228;
  reg [1-1:0] verilogPut_test_1229;
  reg [4-1:0] verilogPut_next_1230;
  reg [4-1:0] verilogPut_root_1231;
  reg [1-1:0] verilogPut_isFree_1232;
  reg [4-1:0] verilogPut_index_1233;
  reg [3-1:0] verilogPut_size_1234;
  reg [1-1:0] verilogPut_isLeaf_1235;
  reg [4-1:0] verilogPut_nextFree_1236;
  reg [64-1:0] verilogPut_Key_0_1237;
  reg [1-1:0] verilogPut_KeyCompares_0_1238;
  reg [3-1:0] verilogPut_KeyCollapse_0_1239;
  reg [8-1:0] verilogPut_Data_0_1240;
  reg [64-1:0] verilogPut_Key_1_1241;
  reg [1-1:0] verilogPut_KeyCompares_1_1242;
  reg [3-1:0] verilogPut_KeyCollapse_1_1243;
  reg [8-1:0] verilogPut_Data_1_1244;
  reg [64-1:0] verilogPut_Key_2_1245;
  reg [1-1:0] verilogPut_KeyCompares_2_1246;
  reg [3-1:0] verilogPut_KeyCollapse_2_1247;
  reg [8-1:0] verilogPut_Data_2_1248;
  reg [64-1:0] verilogPut_Key_3_1249;
  reg [1-1:0] verilogPut_KeyCompares_3_1250;
  reg [3-1:0] verilogPut_KeyCollapse_3_1251;
  reg [8-1:0] verilogPut_Data_3_1252;
  reg [1-1:0] verilogPut_Found_1253;
  reg [64-1:0] verilogPut_Key_1254;
  reg [64-1:0] verilogPut_FoundKey_1255;
  reg [8-1:0] verilogPut_Data_1256;
  reg [4-1:0] verilogPut_BtreeIndex_1257;
  reg [3-1:0] verilogPut_StuckIndex_1258;
  reg [1-1:0] verilogPut_MergeSuccess_1259;
  reg [4-1:0] verilogPut_index_1260;
  reg [3-1:0] verilogPut_size_1261;
  reg [1-1:0] verilogPut_isLeaf_1262;
  reg [4-1:0] verilogPut_nextFree_1263;
  reg [64-1:0] verilogPut_Key_0_1264;
  reg [1-1:0] verilogPut_KeyCompares_0_1265;
  reg [3-1:0] verilogPut_KeyCollapse_0_1266;
  reg [8-1:0] verilogPut_Data_0_1267;
  reg [64-1:0] verilogPut_Key_1_1268;
  reg [1-1:0] verilogPut_KeyCompares_1_1269;
  reg [3-1:0] verilogPut_KeyCollapse_1_1270;
  reg [8-1:0] verilogPut_Data_1_1271;
  reg [64-1:0] verilogPut_Key_2_1272;
  reg [1-1:0] verilogPut_KeyCompares_2_1273;
  reg [3-1:0] verilogPut_KeyCollapse_2_1274;
  reg [8-1:0] verilogPut_Data_2_1275;
  reg [64-1:0] verilogPut_Key_3_1276;
  reg [1-1:0] verilogPut_KeyCompares_3_1277;
  reg [3-1:0] verilogPut_KeyCollapse_3_1278;
  reg [8-1:0] verilogPut_Data_3_1279;
  reg [1-1:0] verilogPut_Found_1280;
  reg [64-1:0] verilogPut_Key_1281;
  reg [64-1:0] verilogPut_FoundKey_1282;
  reg [8-1:0] verilogPut_Data_1283;
  reg [4-1:0] verilogPut_BtreeIndex_1284;
  reg [3-1:0] verilogPut_StuckIndex_1285;
  reg [1-1:0] verilogPut_MergeSuccess_1286;
  reg [64-1:0] verilogPut_childKey_1287;
  reg [4-1:0] verilogPut_childData_1288;
  reg [4-1:0] verilogPut_indexLeft_1289;
  reg [4-1:0] verilogPut_indexRight_1290;
  reg [64-1:0] verilogPut_midKey_1291;
  reg [1-1:0] verilogPut_success_1292;
  reg [1-1:0] verilogPut_test_1293;
  reg [4-1:0] verilogPut_next_1294;
  reg [4-1:0] verilogPut_root_1295;
  reg [1-1:0] verilogPut_isFree_1296;
  reg [4-1:0] verilogPut_index_1297;
  reg [3-1:0] verilogPut_size_1298;
  reg [1-1:0] verilogPut_isLeaf_1299;
  reg [4-1:0] verilogPut_nextFree_1300;
  reg [64-1:0] verilogPut_Key_0_1301;
  reg [1-1:0] verilogPut_KeyCompares_0_1302;
  reg [3-1:0] verilogPut_KeyCollapse_0_1303;
  reg [8-1:0] verilogPut_Data_0_1304;
  reg [64-1:0] verilogPut_Key_1_1305;
  reg [1-1:0] verilogPut_KeyCompares_1_1306;
  reg [3-1:0] verilogPut_KeyCollapse_1_1307;
  reg [8-1:0] verilogPut_Data_1_1308;
  reg [64-1:0] verilogPut_Key_2_1309;
  reg [1-1:0] verilogPut_KeyCompares_2_1310;
  reg [3-1:0] verilogPut_KeyCollapse_2_1311;
  reg [8-1:0] verilogPut_Data_2_1312;
  reg [64-1:0] verilogPut_Key_3_1313;
  reg [1-1:0] verilogPut_KeyCompares_3_1314;
  reg [3-1:0] verilogPut_KeyCollapse_3_1315;
  reg [8-1:0] verilogPut_Data_3_1316;
  reg [1-1:0] verilogPut_Found_1317;
  reg [64-1:0] verilogPut_Key_1318;
  reg [64-1:0] verilogPut_FoundKey_1319;
  reg [8-1:0] verilogPut_Data_1320;
  reg [4-1:0] verilogPut_BtreeIndex_1321;
  reg [3-1:0] verilogPut_StuckIndex_1322;
  reg [1-1:0] verilogPut_MergeSuccess_1323;
  reg [4-1:0] verilogPut_index_1324;
  reg [3-1:0] verilogPut_size_1325;
  reg [1-1:0] verilogPut_isLeaf_1326;
  reg [4-1:0] verilogPut_nextFree_1327;
  reg [64-1:0] verilogPut_Key_0_1328;
  reg [1-1:0] verilogPut_KeyCompares_0_1329;
  reg [3-1:0] verilogPut_KeyCollapse_0_1330;
  reg [8-1:0] verilogPut_Data_0_1331;
  reg [64-1:0] verilogPut_Key_1_1332;
  reg [1-1:0] verilogPut_KeyCompares_1_1333;
  reg [3-1:0] verilogPut_KeyCollapse_1_1334;
  reg [8-1:0] verilogPut_Data_1_1335;
  reg [64-1:0] verilogPut_Key_2_1336;
  reg [1-1:0] verilogPut_KeyCompares_2_1337;
  reg [3-1:0] verilogPut_KeyCollapse_2_1338;
  reg [8-1:0] verilogPut_Data_2_1339;
  reg [64-1:0] verilogPut_Key_3_1340;
  reg [1-1:0] verilogPut_KeyCompares_3_1341;
  reg [3-1:0] verilogPut_KeyCollapse_3_1342;
  reg [8-1:0] verilogPut_Data_3_1343;
  reg [1-1:0] verilogPut_Found_1344;
  reg [64-1:0] verilogPut_Key_1345;
  reg [64-1:0] verilogPut_FoundKey_1346;
  reg [8-1:0] verilogPut_Data_1347;
  reg [4-1:0] verilogPut_BtreeIndex_1348;
  reg [3-1:0] verilogPut_StuckIndex_1349;
  reg [1-1:0] verilogPut_MergeSuccess_1350;
  reg [64-1:0] verilogPut_childKey_1351;
  reg [3-1:0] verilogPut_leftChild_1352;
  reg [3-1:0] verilogPut_rightChild_1353;
  reg [4-1:0] verilogPut_childData_1354;
  reg [4-1:0] verilogPut_indexLeft_1355;
  reg [4-1:0] verilogPut_indexRight_1356;
  reg [64-1:0] verilogPut_midKey_1357;
  reg [1-1:0] verilogPut_success_1358;
  reg [1-1:0] verilogPut_test_1359;
  reg [4-1:0] verilogPut_next_1360;
  reg [4-1:0] verilogPut_root_1361;
  reg [1-1:0] verilogPut_isFree_1362;
  reg [4-1:0] verilogPut_index_1363;
  reg [3-1:0] verilogPut_size_1364;
  reg [1-1:0] verilogPut_isLeaf_1365;
  reg [4-1:0] verilogPut_nextFree_1366;
  reg [64-1:0] verilogPut_Key_0_1367;
  reg [1-1:0] verilogPut_KeyCompares_0_1368;
  reg [3-1:0] verilogPut_KeyCollapse_0_1369;
  reg [8-1:0] verilogPut_Data_0_1370;
  reg [64-1:0] verilogPut_Key_1_1371;
  reg [1-1:0] verilogPut_KeyCompares_1_1372;
  reg [3-1:0] verilogPut_KeyCollapse_1_1373;
  reg [8-1:0] verilogPut_Data_1_1374;
  reg [64-1:0] verilogPut_Key_2_1375;
  reg [1-1:0] verilogPut_KeyCompares_2_1376;
  reg [3-1:0] verilogPut_KeyCollapse_2_1377;
  reg [8-1:0] verilogPut_Data_2_1378;
  reg [64-1:0] verilogPut_Key_3_1379;
  reg [1-1:0] verilogPut_KeyCompares_3_1380;
  reg [3-1:0] verilogPut_KeyCollapse_3_1381;
  reg [8-1:0] verilogPut_Data_3_1382;
  reg [1-1:0] verilogPut_Found_1383;
  reg [64-1:0] verilogPut_Key_1384;
  reg [64-1:0] verilogPut_FoundKey_1385;
  reg [8-1:0] verilogPut_Data_1386;
  reg [4-1:0] verilogPut_BtreeIndex_1387;
  reg [3-1:0] verilogPut_StuckIndex_1388;
  reg [1-1:0] verilogPut_MergeSuccess_1389;
  reg [4-1:0] verilogPut_index_1390;
  reg [3-1:0] verilogPut_size_1391;
  reg [1-1:0] verilogPut_isLeaf_1392;
  reg [4-1:0] verilogPut_nextFree_1393;
  reg [64-1:0] verilogPut_Key_0_1394;
  reg [1-1:0] verilogPut_KeyCompares_0_1395;
  reg [3-1:0] verilogPut_KeyCollapse_0_1396;
  reg [8-1:0] verilogPut_Data_0_1397;
  reg [64-1:0] verilogPut_Key_1_1398;
  reg [1-1:0] verilogPut_KeyCompares_1_1399;
  reg [3-1:0] verilogPut_KeyCollapse_1_1400;
  reg [8-1:0] verilogPut_Data_1_1401;
  reg [64-1:0] verilogPut_Key_2_1402;
  reg [1-1:0] verilogPut_KeyCompares_2_1403;
  reg [3-1:0] verilogPut_KeyCollapse_2_1404;
  reg [8-1:0] verilogPut_Data_2_1405;
  reg [64-1:0] verilogPut_Key_3_1406;
  reg [1-1:0] verilogPut_KeyCompares_3_1407;
  reg [3-1:0] verilogPut_KeyCollapse_3_1408;
  reg [8-1:0] verilogPut_Data_3_1409;
  reg [1-1:0] verilogPut_Found_1410;
  reg [64-1:0] verilogPut_Key_1411;
  reg [64-1:0] verilogPut_FoundKey_1412;
  reg [8-1:0] verilogPut_Data_1413;
  reg [4-1:0] verilogPut_BtreeIndex_1414;
  reg [3-1:0] verilogPut_StuckIndex_1415;
  reg [1-1:0] verilogPut_MergeSuccess_1416;
  reg [64-1:0] verilogPut_childKey_1417;
  reg [4-1:0] verilogPut_childData_1418;
  reg [4-1:0] verilogPut_indexLeft_1419;
  reg [4-1:0] verilogPut_indexRight_1420;
  reg [64-1:0] verilogPut_midKey_1421;
  reg [1-1:0] verilogPut_success_1422;
  reg [1-1:0] verilogPut_test_1423;
  reg [4-1:0] verilogPut_next_1424;
  reg [4-1:0] verilogPut_root_1425;
  reg [1-1:0] verilogPut_isFree_1426;
  reg [4-1:0] verilogPut_index_1427;
  reg [3-1:0] verilogPut_size_1428;
  reg [1-1:0] verilogPut_isLeaf_1429;
  reg [4-1:0] verilogPut_nextFree_1430;
  reg [64-1:0] verilogPut_Key_0_1431;
  reg [1-1:0] verilogPut_KeyCompares_0_1432;
  reg [3-1:0] verilogPut_KeyCollapse_0_1433;
  reg [8-1:0] verilogPut_Data_0_1434;
  reg [64-1:0] verilogPut_Key_1_1435;
  reg [1-1:0] verilogPut_KeyCompares_1_1436;
  reg [3-1:0] verilogPut_KeyCollapse_1_1437;
  reg [8-1:0] verilogPut_Data_1_1438;
  reg [64-1:0] verilogPut_Key_2_1439;
  reg [1-1:0] verilogPut_KeyCompares_2_1440;
  reg [3-1:0] verilogPut_KeyCollapse_2_1441;
  reg [8-1:0] verilogPut_Data_2_1442;
  reg [64-1:0] verilogPut_Key_3_1443;
  reg [1-1:0] verilogPut_KeyCompares_3_1444;
  reg [3-1:0] verilogPut_KeyCollapse_3_1445;
  reg [8-1:0] verilogPut_Data_3_1446;
  reg [1-1:0] verilogPut_Found_1447;
  reg [64-1:0] verilogPut_Key_1448;
  reg [64-1:0] verilogPut_FoundKey_1449;
  reg [8-1:0] verilogPut_Data_1450;
  reg [4-1:0] verilogPut_BtreeIndex_1451;
  reg [3-1:0] verilogPut_StuckIndex_1452;
  reg [1-1:0] verilogPut_MergeSuccess_1453;
  reg [4-1:0] verilogPut_index_1454;
  reg [3-1:0] verilogPut_size_1455;
  reg [1-1:0] verilogPut_isLeaf_1456;
  reg [4-1:0] verilogPut_nextFree_1457;
  reg [64-1:0] verilogPut_Key_0_1458;
  reg [1-1:0] verilogPut_KeyCompares_0_1459;
  reg [3-1:0] verilogPut_KeyCollapse_0_1460;
  reg [8-1:0] verilogPut_Data_0_1461;
  reg [64-1:0] verilogPut_Key_1_1462;
  reg [1-1:0] verilogPut_KeyCompares_1_1463;
  reg [3-1:0] verilogPut_KeyCollapse_1_1464;
  reg [8-1:0] verilogPut_Data_1_1465;
  reg [64-1:0] verilogPut_Key_2_1466;
  reg [1-1:0] verilogPut_KeyCompares_2_1467;
  reg [3-1:0] verilogPut_KeyCollapse_2_1468;
  reg [8-1:0] verilogPut_Data_2_1469;
  reg [64-1:0] verilogPut_Key_3_1470;
  reg [1-1:0] verilogPut_KeyCompares_3_1471;
  reg [3-1:0] verilogPut_KeyCollapse_3_1472;
  reg [8-1:0] verilogPut_Data_3_1473;
  reg [1-1:0] verilogPut_Found_1474;
  reg [64-1:0] verilogPut_Key_1475;
  reg [64-1:0] verilogPut_FoundKey_1476;
  reg [8-1:0] verilogPut_Data_1477;
  reg [4-1:0] verilogPut_BtreeIndex_1478;
  reg [3-1:0] verilogPut_StuckIndex_1479;
  reg [1-1:0] verilogPut_MergeSuccess_1480;
  reg [64-1:0] verilogPut_childKey_1481;
  reg [3-1:0] verilogPut_leftChild_1482;
  reg [3-1:0] verilogPut_rightChild_1483;
  reg [4-1:0] verilogPut_childData_1484;
  reg [4-1:0] verilogPut_indexLeft_1485;
  reg [4-1:0] verilogPut_indexRight_1486;
  reg [64-1:0] verilogPut_midKey_1487;
  reg [1-1:0] verilogPut_success_1488;
  reg [1-1:0] verilogPut_test_1489;
  reg [4-1:0] verilogPut_next_1490;
  reg [4-1:0] verilogPut_root_1491;
  reg [1-1:0] verilogPut_isFree_1492;
  integer verilogPut_pc;
  integer verilogPut_stop;
  integer verilogPut_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      verilogPut_pc <= 0;
      verilogPut_stop <= 0;
      verilogPut_returnCode <= 0;
      verilogPut_index_2 <= 0;
      verilogPut_size_3 <= 0;
      verilogPut_isLeaf_4 <= 0;
      verilogPut_nextFree_5 <= 0;
      verilogPut_Key_0_6 <= 0;
      verilogPut_KeyCompares_0_7 <= 0;
      verilogPut_KeyCollapse_0_8 <= 0;
      verilogPut_Data_0_9 <= 0;
      verilogPut_stuckKeys_0_1_index_10 <= 0;
      verilogPut_stuckKeys_0_2_index_11 <= 0;
      verilogPut_stuckKeys_0_2_value_12 <= 0;
      verilogPut_stuckData_0_3_index_13 <= 0;
      verilogPut_stuckData_0_4_index_14 <= 0;
      verilogPut_stuckData_0_4_value_15 <= 0;
      verilogPut_Key_1_16 <= 0;
      verilogPut_KeyCompares_1_17 <= 0;
      verilogPut_KeyCollapse_1_18 <= 0;
      verilogPut_Data_1_19 <= 0;
      verilogPut_stuckKeys_1_5_index_20 <= 0;
      verilogPut_stuckKeys_1_6_index_21 <= 0;
      verilogPut_stuckKeys_1_6_value_22 <= 0;
      verilogPut_stuckData_1_7_index_23 <= 0;
      verilogPut_stuckData_1_8_index_24 <= 0;
      verilogPut_stuckData_1_8_value_25 <= 0;
      verilogPut_Key_2_26 <= 0;
      verilogPut_KeyCompares_2_27 <= 0;
      verilogPut_KeyCollapse_2_28 <= 0;
      verilogPut_Data_2_29 <= 0;
      verilogPut_stuckKeys_2_9_index_30 <= 0;
      verilogPut_stuckKeys_2_10_index_31 <= 0;
      verilogPut_stuckKeys_2_10_value_32 <= 0;
      verilogPut_stuckData_2_11_index_33 <= 0;
      verilogPut_stuckData_2_12_index_34 <= 0;
      verilogPut_stuckData_2_12_value_35 <= 0;
      verilogPut_Key_3_36 <= 0;
      verilogPut_KeyCompares_3_37 <= 0;
      verilogPut_KeyCollapse_3_38 <= 0;
      verilogPut_Data_3_39 <= 0;
      verilogPut_stuckKeys_3_13_index_40 <= 0;
      verilogPut_stuckKeys_3_14_index_41 <= 0;
      verilogPut_stuckKeys_3_14_value_42 <= 0;
      verilogPut_stuckData_3_15_index_43 <= 0;
      verilogPut_stuckData_3_16_index_44 <= 0;
      verilogPut_stuckData_3_16_value_45 <= 0;
      verilogPut_stuckSize_17_index_46 <= 0;
      verilogPut_stuckSize_18_index_47 <= 0;
      verilogPut_stuckSize_18_value_48 <= 0;
      verilogPut_stuckIsLeaf_19_index_49 <= 0;
      verilogPut_stuckIsLeaf_20_index_50 <= 0;
      verilogPut_stuckIsLeaf_20_value_51 <= 0;
      verilogPut_Found_52 <= 0;
      verilogPut_Key_53 <= 0;
      verilogPut_FoundKey_54 <= 0;
      verilogPut_Data_55 <= 0;
      verilogPut_BtreeIndex_56 <= 0;
      verilogPut_StuckIndex_57 <= 0;
      verilogPut_MergeSuccess_58 <= 0;
      verilogPut_index_59 <= 0;
      verilogPut_size_60 <= 0;
      verilogPut_isLeaf_61 <= 0;
      verilogPut_nextFree_62 <= 0;
      verilogPut_Key_0_63 <= 0;
      verilogPut_KeyCompares_0_64 <= 0;
      verilogPut_KeyCollapse_0_65 <= 0;
      verilogPut_Data_0_66 <= 0;
      verilogPut_Key_1_67 <= 0;
      verilogPut_KeyCompares_1_68 <= 0;
      verilogPut_KeyCollapse_1_69 <= 0;
      verilogPut_Data_1_70 <= 0;
      verilogPut_Key_2_71 <= 0;
      verilogPut_KeyCompares_2_72 <= 0;
      verilogPut_KeyCollapse_2_73 <= 0;
      verilogPut_Data_2_74 <= 0;
      verilogPut_Key_3_75 <= 0;
      verilogPut_KeyCompares_3_76 <= 0;
      verilogPut_KeyCollapse_3_77 <= 0;
      verilogPut_Data_3_78 <= 0;
      verilogPut_Found_79 <= 0;
      verilogPut_Key_80 <= 0;
      verilogPut_FoundKey_81 <= 0;
      verilogPut_Data_82 <= 0;
      verilogPut_BtreeIndex_83 <= 0;
      verilogPut_StuckIndex_84 <= 0;
      verilogPut_MergeSuccess_85 <= 0;
      verilogPut_index_86 <= 0;
      verilogPut_size_87 <= 0;
      verilogPut_isLeaf_88 <= 0;
      verilogPut_nextFree_89 <= 0;
      verilogPut_Key_0_90 <= 0;
      verilogPut_KeyCompares_0_91 <= 0;
      verilogPut_KeyCollapse_0_92 <= 0;
      verilogPut_Data_0_93 <= 0;
      verilogPut_Key_1_94 <= 0;
      verilogPut_KeyCompares_1_95 <= 0;
      verilogPut_KeyCollapse_1_96 <= 0;
      verilogPut_Data_1_97 <= 0;
      verilogPut_Key_2_98 <= 0;
      verilogPut_KeyCompares_2_99 <= 0;
      verilogPut_KeyCollapse_2_100 <= 0;
      verilogPut_Data_2_101 <= 0;
      verilogPut_Key_3_102 <= 0;
      verilogPut_KeyCompares_3_103 <= 0;
      verilogPut_KeyCollapse_3_104 <= 0;
      verilogPut_Data_3_105 <= 0;
      verilogPut_Found_106 <= 0;
      verilogPut_Key_107 <= 0;
      verilogPut_FoundKey_108 <= 0;
      verilogPut_Data_109 <= 0;
      verilogPut_BtreeIndex_110 <= 0;
      verilogPut_StuckIndex_111 <= 0;
      verilogPut_MergeSuccess_112 <= 0;
      verilogPut_child_113 <= 0;
      verilogPut_parent_114 <= 0;
      verilogPut_childInparent_115 <= 0;
      verilogPut_found_116 <= 0;
      verilogPut_full_117 <= 0;
      verilogPut_i_118 <= 0;
      verilogPut_notFull_119 <= 0;
      verilogPut_index_120 <= 0;
      verilogPut_size_121 <= 0;
      verilogPut_isLeaf_122 <= 0;
      verilogPut_nextFree_123 <= 0;
      verilogPut_Key_0_124 <= 0;
      verilogPut_KeyCompares_0_125 <= 0;
      verilogPut_KeyCollapse_0_126 <= 0;
      verilogPut_Data_0_127 <= 0;
      verilogPut_Key_1_128 <= 0;
      verilogPut_KeyCompares_1_129 <= 0;
      verilogPut_KeyCollapse_1_130 <= 0;
      verilogPut_Data_1_131 <= 0;
      verilogPut_Key_2_132 <= 0;
      verilogPut_KeyCompares_2_133 <= 0;
      verilogPut_KeyCollapse_2_134 <= 0;
      verilogPut_Data_2_135 <= 0;
      verilogPut_Key_3_136 <= 0;
      verilogPut_KeyCompares_3_137 <= 0;
      verilogPut_KeyCollapse_3_138 <= 0;
      verilogPut_Data_3_139 <= 0;
      verilogPut_Found_140 <= 0;
      verilogPut_Key_141 <= 0;
      verilogPut_FoundKey_142 <= 0;
      verilogPut_Data_143 <= 0;
      verilogPut_BtreeIndex_144 <= 0;
      verilogPut_StuckIndex_145 <= 0;
      verilogPut_MergeSuccess_146 <= 0;
      verilogPut_index_147 <= 0;
      verilogPut_size_148 <= 0;
      verilogPut_isLeaf_149 <= 0;
      verilogPut_nextFree_150 <= 0;
      verilogPut_Key_0_151 <= 0;
      verilogPut_KeyCompares_0_152 <= 0;
      verilogPut_KeyCollapse_0_153 <= 0;
      verilogPut_Data_0_154 <= 0;
      verilogPut_Key_1_155 <= 0;
      verilogPut_KeyCompares_1_156 <= 0;
      verilogPut_KeyCollapse_1_157 <= 0;
      verilogPut_Data_1_158 <= 0;
      verilogPut_Key_2_159 <= 0;
      verilogPut_KeyCompares_2_160 <= 0;
      verilogPut_KeyCollapse_2_161 <= 0;
      verilogPut_Data_2_162 <= 0;
      verilogPut_Key_3_163 <= 0;
      verilogPut_KeyCompares_3_164 <= 0;
      verilogPut_KeyCollapse_3_165 <= 0;
      verilogPut_Data_3_166 <= 0;
      verilogPut_Found_167 <= 0;
      verilogPut_Key_168 <= 0;
      verilogPut_FoundKey_169 <= 0;
      verilogPut_Data_170 <= 0;
      verilogPut_BtreeIndex_171 <= 0;
      verilogPut_StuckIndex_172 <= 0;
      verilogPut_MergeSuccess_173 <= 0;
      verilogPut_index_174 <= 0;
      verilogPut_size_175 <= 0;
      verilogPut_isLeaf_176 <= 0;
      verilogPut_nextFree_177 <= 0;
      verilogPut_Key_0_178 <= 0;
      verilogPut_KeyCompares_0_179 <= 0;
      verilogPut_KeyCollapse_0_180 <= 0;
      verilogPut_Data_0_181 <= 0;
      verilogPut_Key_1_182 <= 0;
      verilogPut_KeyCompares_1_183 <= 0;
      verilogPut_KeyCollapse_1_184 <= 0;
      verilogPut_Data_1_185 <= 0;
      verilogPut_Key_2_186 <= 0;
      verilogPut_KeyCompares_2_187 <= 0;
      verilogPut_KeyCollapse_2_188 <= 0;
      verilogPut_Data_2_189 <= 0;
      verilogPut_Key_3_190 <= 0;
      verilogPut_KeyCompares_3_191 <= 0;
      verilogPut_KeyCollapse_3_192 <= 0;
      verilogPut_Data_3_193 <= 0;
      verilogPut_Found_194 <= 0;
      verilogPut_Key_195 <= 0;
      verilogPut_FoundKey_196 <= 0;
      verilogPut_Data_197 <= 0;
      verilogPut_BtreeIndex_198 <= 0;
      verilogPut_StuckIndex_199 <= 0;
      verilogPut_MergeSuccess_200 <= 0;
      verilogPut_indexLeft_201 <= 0;
      verilogPut_indexRight_202 <= 0;
      verilogPut_midKey_203 <= 0;
      verilogPut_freeNext_21_index_204 <= 0;
      verilogPut_freeNext_22_index_205 <= 0;
      verilogPut_freeNext_22_value_206 <= 0;
      verilogPut_stuckIsFree_23_index_207 <= 0;
      verilogPut_stuckIsFree_23_value_208 <= 0;
      verilogPut_root_209 <= 0;
      verilogPut_next_210 <= 0;
      verilogPut_isLeaf_211 <= 0;
      verilogPut_isFree_212 <= 0;
      verilogPut_root_213 <= 0;
      verilogPut_next_214 <= 0;
      verilogPut_isLeaf_215 <= 0;
      verilogPut_isFree_216 <= 0;
      verilogPut_i_217 <= 0;
      verilogPut_notFull_218 <= 0;
      verilogPut_index_219 <= 0;
      verilogPut_size_220 <= 0;
      verilogPut_isLeaf_221 <= 0;
      verilogPut_nextFree_222 <= 0;
      verilogPut_Key_0_223 <= 0;
      verilogPut_KeyCompares_0_224 <= 0;
      verilogPut_KeyCollapse_0_225 <= 0;
      verilogPut_Data_0_226 <= 0;
      verilogPut_Key_1_227 <= 0;
      verilogPut_KeyCompares_1_228 <= 0;
      verilogPut_KeyCollapse_1_229 <= 0;
      verilogPut_Data_1_230 <= 0;
      verilogPut_Key_2_231 <= 0;
      verilogPut_KeyCompares_2_232 <= 0;
      verilogPut_KeyCollapse_2_233 <= 0;
      verilogPut_Data_2_234 <= 0;
      verilogPut_Key_3_235 <= 0;
      verilogPut_KeyCompares_3_236 <= 0;
      verilogPut_KeyCollapse_3_237 <= 0;
      verilogPut_Data_3_238 <= 0;
      verilogPut_Found_239 <= 0;
      verilogPut_Key_240 <= 0;
      verilogPut_FoundKey_241 <= 0;
      verilogPut_Data_242 <= 0;
      verilogPut_BtreeIndex_243 <= 0;
      verilogPut_StuckIndex_244 <= 0;
      verilogPut_MergeSuccess_245 <= 0;
      verilogPut_index_246 <= 0;
      verilogPut_size_247 <= 0;
      verilogPut_isLeaf_248 <= 0;
      verilogPut_nextFree_249 <= 0;
      verilogPut_Key_0_250 <= 0;
      verilogPut_KeyCompares_0_251 <= 0;
      verilogPut_KeyCollapse_0_252 <= 0;
      verilogPut_Data_0_253 <= 0;
      verilogPut_Key_1_254 <= 0;
      verilogPut_KeyCompares_1_255 <= 0;
      verilogPut_KeyCollapse_1_256 <= 0;
      verilogPut_Data_1_257 <= 0;
      verilogPut_Key_2_258 <= 0;
      verilogPut_KeyCompares_2_259 <= 0;
      verilogPut_KeyCollapse_2_260 <= 0;
      verilogPut_Data_2_261 <= 0;
      verilogPut_Key_3_262 <= 0;
      verilogPut_KeyCompares_3_263 <= 0;
      verilogPut_KeyCollapse_3_264 <= 0;
      verilogPut_Data_3_265 <= 0;
      verilogPut_Found_266 <= 0;
      verilogPut_Key_267 <= 0;
      verilogPut_FoundKey_268 <= 0;
      verilogPut_Data_269 <= 0;
      verilogPut_BtreeIndex_270 <= 0;
      verilogPut_StuckIndex_271 <= 0;
      verilogPut_MergeSuccess_272 <= 0;
      verilogPut_index_273 <= 0;
      verilogPut_size_274 <= 0;
      verilogPut_isLeaf_275 <= 0;
      verilogPut_nextFree_276 <= 0;
      verilogPut_Key_0_277 <= 0;
      verilogPut_KeyCompares_0_278 <= 0;
      verilogPut_KeyCollapse_0_279 <= 0;
      verilogPut_Data_0_280 <= 0;
      verilogPut_Key_1_281 <= 0;
      verilogPut_KeyCompares_1_282 <= 0;
      verilogPut_KeyCollapse_1_283 <= 0;
      verilogPut_Data_1_284 <= 0;
      verilogPut_Key_2_285 <= 0;
      verilogPut_KeyCompares_2_286 <= 0;
      verilogPut_KeyCollapse_2_287 <= 0;
      verilogPut_Data_2_288 <= 0;
      verilogPut_Key_3_289 <= 0;
      verilogPut_KeyCompares_3_290 <= 0;
      verilogPut_KeyCollapse_3_291 <= 0;
      verilogPut_Data_3_292 <= 0;
      verilogPut_Found_293 <= 0;
      verilogPut_Key_294 <= 0;
      verilogPut_FoundKey_295 <= 0;
      verilogPut_Data_296 <= 0;
      verilogPut_BtreeIndex_297 <= 0;
      verilogPut_StuckIndex_298 <= 0;
      verilogPut_MergeSuccess_299 <= 0;
      verilogPut_indexLeft_300 <= 0;
      verilogPut_indexRight_301 <= 0;
      verilogPut_midKey_302 <= 0;
      verilogPut_root_303 <= 0;
      verilogPut_next_304 <= 0;
      verilogPut_isLeaf_305 <= 0;
      verilogPut_isFree_306 <= 0;
      verilogPut_root_307 <= 0;
      verilogPut_next_308 <= 0;
      verilogPut_isLeaf_309 <= 0;
      verilogPut_isFree_310 <= 0;
      verilogPut_index_311 <= 0;
      verilogPut_size_312 <= 0;
      verilogPut_isLeaf_313 <= 0;
      verilogPut_nextFree_314 <= 0;
      verilogPut_Key_0_315 <= 0;
      verilogPut_KeyCompares_0_316 <= 0;
      verilogPut_KeyCollapse_0_317 <= 0;
      verilogPut_Data_0_318 <= 0;
      verilogPut_Key_1_319 <= 0;
      verilogPut_KeyCompares_1_320 <= 0;
      verilogPut_KeyCollapse_1_321 <= 0;
      verilogPut_Data_1_322 <= 0;
      verilogPut_Key_2_323 <= 0;
      verilogPut_KeyCompares_2_324 <= 0;
      verilogPut_KeyCollapse_2_325 <= 0;
      verilogPut_Data_2_326 <= 0;
      verilogPut_Key_3_327 <= 0;
      verilogPut_KeyCompares_3_328 <= 0;
      verilogPut_KeyCollapse_3_329 <= 0;
      verilogPut_Data_3_330 <= 0;
      verilogPut_Found_331 <= 0;
      verilogPut_Key_332 <= 0;
      verilogPut_FoundKey_333 <= 0;
      verilogPut_Data_334 <= 0;
      verilogPut_BtreeIndex_335 <= 0;
      verilogPut_StuckIndex_336 <= 0;
      verilogPut_MergeSuccess_337 <= 0;
      verilogPut_index_338 <= 0;
      verilogPut_size_339 <= 0;
      verilogPut_isLeaf_340 <= 0;
      verilogPut_nextFree_341 <= 0;
      verilogPut_Key_0_342 <= 0;
      verilogPut_KeyCompares_0_343 <= 0;
      verilogPut_KeyCollapse_0_344 <= 0;
      verilogPut_Data_0_345 <= 0;
      verilogPut_Key_1_346 <= 0;
      verilogPut_KeyCompares_1_347 <= 0;
      verilogPut_KeyCollapse_1_348 <= 0;
      verilogPut_Data_1_349 <= 0;
      verilogPut_Key_2_350 <= 0;
      verilogPut_KeyCompares_2_351 <= 0;
      verilogPut_KeyCollapse_2_352 <= 0;
      verilogPut_Data_2_353 <= 0;
      verilogPut_Key_3_354 <= 0;
      verilogPut_KeyCompares_3_355 <= 0;
      verilogPut_KeyCollapse_3_356 <= 0;
      verilogPut_Data_3_357 <= 0;
      verilogPut_Found_358 <= 0;
      verilogPut_Key_359 <= 0;
      verilogPut_FoundKey_360 <= 0;
      verilogPut_Data_361 <= 0;
      verilogPut_BtreeIndex_362 <= 0;
      verilogPut_StuckIndex_363 <= 0;
      verilogPut_MergeSuccess_364 <= 0;
      verilogPut_index_365 <= 0;
      verilogPut_size_366 <= 0;
      verilogPut_isLeaf_367 <= 0;
      verilogPut_nextFree_368 <= 0;
      verilogPut_Key_0_369 <= 0;
      verilogPut_KeyCompares_0_370 <= 0;
      verilogPut_KeyCollapse_0_371 <= 0;
      verilogPut_Data_0_372 <= 0;
      verilogPut_Key_1_373 <= 0;
      verilogPut_KeyCompares_1_374 <= 0;
      verilogPut_KeyCollapse_1_375 <= 0;
      verilogPut_Data_1_376 <= 0;
      verilogPut_Key_2_377 <= 0;
      verilogPut_KeyCompares_2_378 <= 0;
      verilogPut_KeyCollapse_2_379 <= 0;
      verilogPut_Data_2_380 <= 0;
      verilogPut_Key_3_381 <= 0;
      verilogPut_KeyCompares_3_382 <= 0;
      verilogPut_KeyCollapse_3_383 <= 0;
      verilogPut_Data_3_384 <= 0;
      verilogPut_Found_385 <= 0;
      verilogPut_Key_386 <= 0;
      verilogPut_FoundKey_387 <= 0;
      verilogPut_Data_388 <= 0;
      verilogPut_BtreeIndex_389 <= 0;
      verilogPut_StuckIndex_390 <= 0;
      verilogPut_MergeSuccess_391 <= 0;
      verilogPut_index_392 <= 0;
      verilogPut_size_393 <= 0;
      verilogPut_isLeaf_394 <= 0;
      verilogPut_nextFree_395 <= 0;
      verilogPut_Key_0_396 <= 0;
      verilogPut_KeyCompares_0_397 <= 0;
      verilogPut_KeyCollapse_0_398 <= 0;
      verilogPut_Data_0_399 <= 0;
      verilogPut_Key_1_400 <= 0;
      verilogPut_KeyCompares_1_401 <= 0;
      verilogPut_KeyCollapse_1_402 <= 0;
      verilogPut_Data_1_403 <= 0;
      verilogPut_Key_2_404 <= 0;
      verilogPut_KeyCompares_2_405 <= 0;
      verilogPut_KeyCollapse_2_406 <= 0;
      verilogPut_Data_2_407 <= 0;
      verilogPut_Key_3_408 <= 0;
      verilogPut_KeyCompares_3_409 <= 0;
      verilogPut_KeyCollapse_3_410 <= 0;
      verilogPut_Data_3_411 <= 0;
      verilogPut_Found_412 <= 0;
      verilogPut_Key_413 <= 0;
      verilogPut_FoundKey_414 <= 0;
      verilogPut_Data_415 <= 0;
      verilogPut_BtreeIndex_416 <= 0;
      verilogPut_StuckIndex_417 <= 0;
      verilogPut_MergeSuccess_418 <= 0;
      verilogPut_childKey_419 <= 0;
      verilogPut_childData_420 <= 0;
      verilogPut_indexLeft_421 <= 0;
      verilogPut_indexRight_422 <= 0;
      verilogPut_midKey_423 <= 0;
      verilogPut_root_424 <= 0;
      verilogPut_next_425 <= 0;
      verilogPut_isLeaf_426 <= 0;
      verilogPut_isFree_427 <= 0;
      verilogPut_index_428 <= 0;
      verilogPut_size_429 <= 0;
      verilogPut_isLeaf_430 <= 0;
      verilogPut_nextFree_431 <= 0;
      verilogPut_Key_0_432 <= 0;
      verilogPut_KeyCompares_0_433 <= 0;
      verilogPut_KeyCollapse_0_434 <= 0;
      verilogPut_Data_0_435 <= 0;
      verilogPut_Key_1_436 <= 0;
      verilogPut_KeyCompares_1_437 <= 0;
      verilogPut_KeyCollapse_1_438 <= 0;
      verilogPut_Data_1_439 <= 0;
      verilogPut_Key_2_440 <= 0;
      verilogPut_KeyCompares_2_441 <= 0;
      verilogPut_KeyCollapse_2_442 <= 0;
      verilogPut_Data_2_443 <= 0;
      verilogPut_Key_3_444 <= 0;
      verilogPut_KeyCompares_3_445 <= 0;
      verilogPut_KeyCollapse_3_446 <= 0;
      verilogPut_Data_3_447 <= 0;
      verilogPut_Found_448 <= 0;
      verilogPut_Key_449 <= 0;
      verilogPut_FoundKey_450 <= 0;
      verilogPut_Data_451 <= 0;
      verilogPut_BtreeIndex_452 <= 0;
      verilogPut_StuckIndex_453 <= 0;
      verilogPut_MergeSuccess_454 <= 0;
      verilogPut_index_455 <= 0;
      verilogPut_size_456 <= 0;
      verilogPut_isLeaf_457 <= 0;
      verilogPut_nextFree_458 <= 0;
      verilogPut_Key_0_459 <= 0;
      verilogPut_KeyCompares_0_460 <= 0;
      verilogPut_KeyCollapse_0_461 <= 0;
      verilogPut_Data_0_462 <= 0;
      verilogPut_Key_1_463 <= 0;
      verilogPut_KeyCompares_1_464 <= 0;
      verilogPut_KeyCollapse_1_465 <= 0;
      verilogPut_Data_1_466 <= 0;
      verilogPut_Key_2_467 <= 0;
      verilogPut_KeyCompares_2_468 <= 0;
      verilogPut_KeyCollapse_2_469 <= 0;
      verilogPut_Data_2_470 <= 0;
      verilogPut_Key_3_471 <= 0;
      verilogPut_KeyCompares_3_472 <= 0;
      verilogPut_KeyCollapse_3_473 <= 0;
      verilogPut_Data_3_474 <= 0;
      verilogPut_Found_475 <= 0;
      verilogPut_Key_476 <= 0;
      verilogPut_FoundKey_477 <= 0;
      verilogPut_Data_478 <= 0;
      verilogPut_BtreeIndex_479 <= 0;
      verilogPut_StuckIndex_480 <= 0;
      verilogPut_MergeSuccess_481 <= 0;
      verilogPut_index_482 <= 0;
      verilogPut_size_483 <= 0;
      verilogPut_isLeaf_484 <= 0;
      verilogPut_nextFree_485 <= 0;
      verilogPut_Key_0_486 <= 0;
      verilogPut_KeyCompares_0_487 <= 0;
      verilogPut_KeyCollapse_0_488 <= 0;
      verilogPut_Data_0_489 <= 0;
      verilogPut_Key_1_490 <= 0;
      verilogPut_KeyCompares_1_491 <= 0;
      verilogPut_KeyCollapse_1_492 <= 0;
      verilogPut_Data_1_493 <= 0;
      verilogPut_Key_2_494 <= 0;
      verilogPut_KeyCompares_2_495 <= 0;
      verilogPut_KeyCollapse_2_496 <= 0;
      verilogPut_Data_2_497 <= 0;
      verilogPut_Key_3_498 <= 0;
      verilogPut_KeyCompares_3_499 <= 0;
      verilogPut_KeyCollapse_3_500 <= 0;
      verilogPut_Data_3_501 <= 0;
      verilogPut_Found_502 <= 0;
      verilogPut_Key_503 <= 0;
      verilogPut_FoundKey_504 <= 0;
      verilogPut_Data_505 <= 0;
      verilogPut_BtreeIndex_506 <= 0;
      verilogPut_StuckIndex_507 <= 0;
      verilogPut_MergeSuccess_508 <= 0;
      verilogPut_childIndex_509 <= 0;
      verilogPut_leftIndex_510 <= 0;
      verilogPut_midKey_511 <= 0;
      verilogPut_root_512 <= 0;
      verilogPut_next_513 <= 0;
      verilogPut_isLeaf_514 <= 0;
      verilogPut_isFree_515 <= 0;
      verilogPut_i_516 <= 0;
      verilogPut_notFull_517 <= 0;
      verilogPut_index_518 <= 0;
      verilogPut_size_519 <= 0;
      verilogPut_isLeaf_520 <= 0;
      verilogPut_nextFree_521 <= 0;
      verilogPut_Key_0_522 <= 0;
      verilogPut_KeyCompares_0_523 <= 0;
      verilogPut_KeyCollapse_0_524 <= 0;
      verilogPut_Data_0_525 <= 0;
      verilogPut_Key_1_526 <= 0;
      verilogPut_KeyCompares_1_527 <= 0;
      verilogPut_KeyCollapse_1_528 <= 0;
      verilogPut_Data_1_529 <= 0;
      verilogPut_Key_2_530 <= 0;
      verilogPut_KeyCompares_2_531 <= 0;
      verilogPut_KeyCollapse_2_532 <= 0;
      verilogPut_Data_2_533 <= 0;
      verilogPut_Key_3_534 <= 0;
      verilogPut_KeyCompares_3_535 <= 0;
      verilogPut_KeyCollapse_3_536 <= 0;
      verilogPut_Data_3_537 <= 0;
      verilogPut_Found_538 <= 0;
      verilogPut_Key_539 <= 0;
      verilogPut_FoundKey_540 <= 0;
      verilogPut_Data_541 <= 0;
      verilogPut_BtreeIndex_542 <= 0;
      verilogPut_StuckIndex_543 <= 0;
      verilogPut_MergeSuccess_544 <= 0;
      verilogPut_index_545 <= 0;
      verilogPut_size_546 <= 0;
      verilogPut_isLeaf_547 <= 0;
      verilogPut_nextFree_548 <= 0;
      verilogPut_Key_0_549 <= 0;
      verilogPut_KeyCompares_0_550 <= 0;
      verilogPut_KeyCollapse_0_551 <= 0;
      verilogPut_Data_0_552 <= 0;
      verilogPut_Key_1_553 <= 0;
      verilogPut_KeyCompares_1_554 <= 0;
      verilogPut_KeyCollapse_1_555 <= 0;
      verilogPut_Data_1_556 <= 0;
      verilogPut_Key_2_557 <= 0;
      verilogPut_KeyCompares_2_558 <= 0;
      verilogPut_KeyCollapse_2_559 <= 0;
      verilogPut_Data_2_560 <= 0;
      verilogPut_Key_3_561 <= 0;
      verilogPut_KeyCompares_3_562 <= 0;
      verilogPut_KeyCollapse_3_563 <= 0;
      verilogPut_Data_3_564 <= 0;
      verilogPut_Found_565 <= 0;
      verilogPut_Key_566 <= 0;
      verilogPut_FoundKey_567 <= 0;
      verilogPut_Data_568 <= 0;
      verilogPut_BtreeIndex_569 <= 0;
      verilogPut_StuckIndex_570 <= 0;
      verilogPut_MergeSuccess_571 <= 0;
      verilogPut_index_572 <= 0;
      verilogPut_size_573 <= 0;
      verilogPut_isLeaf_574 <= 0;
      verilogPut_nextFree_575 <= 0;
      verilogPut_Key_0_576 <= 0;
      verilogPut_KeyCompares_0_577 <= 0;
      verilogPut_KeyCollapse_0_578 <= 0;
      verilogPut_Data_0_579 <= 0;
      verilogPut_Key_1_580 <= 0;
      verilogPut_KeyCompares_1_581 <= 0;
      verilogPut_KeyCollapse_1_582 <= 0;
      verilogPut_Data_1_583 <= 0;
      verilogPut_Key_2_584 <= 0;
      verilogPut_KeyCompares_2_585 <= 0;
      verilogPut_KeyCollapse_2_586 <= 0;
      verilogPut_Data_2_587 <= 0;
      verilogPut_Key_3_588 <= 0;
      verilogPut_KeyCompares_3_589 <= 0;
      verilogPut_KeyCollapse_3_590 <= 0;
      verilogPut_Data_3_591 <= 0;
      verilogPut_Found_592 <= 0;
      verilogPut_Key_593 <= 0;
      verilogPut_FoundKey_594 <= 0;
      verilogPut_Data_595 <= 0;
      verilogPut_BtreeIndex_596 <= 0;
      verilogPut_StuckIndex_597 <= 0;
      verilogPut_MergeSuccess_598 <= 0;
      verilogPut_index_599 <= 0;
      verilogPut_size_600 <= 0;
      verilogPut_isLeaf_601 <= 0;
      verilogPut_nextFree_602 <= 0;
      verilogPut_Key_0_603 <= 0;
      verilogPut_KeyCompares_0_604 <= 0;
      verilogPut_KeyCollapse_0_605 <= 0;
      verilogPut_Data_0_606 <= 0;
      verilogPut_Key_1_607 <= 0;
      verilogPut_KeyCompares_1_608 <= 0;
      verilogPut_KeyCollapse_1_609 <= 0;
      verilogPut_Data_1_610 <= 0;
      verilogPut_Key_2_611 <= 0;
      verilogPut_KeyCompares_2_612 <= 0;
      verilogPut_KeyCollapse_2_613 <= 0;
      verilogPut_Data_2_614 <= 0;
      verilogPut_Key_3_615 <= 0;
      verilogPut_KeyCompares_3_616 <= 0;
      verilogPut_KeyCollapse_3_617 <= 0;
      verilogPut_Data_3_618 <= 0;
      verilogPut_Found_619 <= 0;
      verilogPut_Key_620 <= 0;
      verilogPut_FoundKey_621 <= 0;
      verilogPut_Data_622 <= 0;
      verilogPut_BtreeIndex_623 <= 0;
      verilogPut_StuckIndex_624 <= 0;
      verilogPut_MergeSuccess_625 <= 0;
      verilogPut_childKey_626 <= 0;
      verilogPut_childData_627 <= 0;
      verilogPut_indexLeft_628 <= 0;
      verilogPut_indexRight_629 <= 0;
      verilogPut_midKey_630 <= 0;
      verilogPut_root_631 <= 0;
      verilogPut_next_632 <= 0;
      verilogPut_isLeaf_633 <= 0;
      verilogPut_isFree_634 <= 0;
      verilogPut_index_635 <= 0;
      verilogPut_size_636 <= 0;
      verilogPut_isLeaf_637 <= 0;
      verilogPut_nextFree_638 <= 0;
      verilogPut_Key_0_639 <= 0;
      verilogPut_KeyCompares_0_640 <= 0;
      verilogPut_KeyCollapse_0_641 <= 0;
      verilogPut_Data_0_642 <= 0;
      verilogPut_Key_1_643 <= 0;
      verilogPut_KeyCompares_1_644 <= 0;
      verilogPut_KeyCollapse_1_645 <= 0;
      verilogPut_Data_1_646 <= 0;
      verilogPut_Key_2_647 <= 0;
      verilogPut_KeyCompares_2_648 <= 0;
      verilogPut_KeyCollapse_2_649 <= 0;
      verilogPut_Data_2_650 <= 0;
      verilogPut_Key_3_651 <= 0;
      verilogPut_KeyCompares_3_652 <= 0;
      verilogPut_KeyCollapse_3_653 <= 0;
      verilogPut_Data_3_654 <= 0;
      verilogPut_Found_655 <= 0;
      verilogPut_Key_656 <= 0;
      verilogPut_FoundKey_657 <= 0;
      verilogPut_Data_658 <= 0;
      verilogPut_BtreeIndex_659 <= 0;
      verilogPut_StuckIndex_660 <= 0;
      verilogPut_MergeSuccess_661 <= 0;
      verilogPut_index_662 <= 0;
      verilogPut_size_663 <= 0;
      verilogPut_isLeaf_664 <= 0;
      verilogPut_nextFree_665 <= 0;
      verilogPut_Key_0_666 <= 0;
      verilogPut_KeyCompares_0_667 <= 0;
      verilogPut_KeyCollapse_0_668 <= 0;
      verilogPut_Data_0_669 <= 0;
      verilogPut_Key_1_670 <= 0;
      verilogPut_KeyCompares_1_671 <= 0;
      verilogPut_KeyCollapse_1_672 <= 0;
      verilogPut_Data_1_673 <= 0;
      verilogPut_Key_2_674 <= 0;
      verilogPut_KeyCompares_2_675 <= 0;
      verilogPut_KeyCollapse_2_676 <= 0;
      verilogPut_Data_2_677 <= 0;
      verilogPut_Key_3_678 <= 0;
      verilogPut_KeyCompares_3_679 <= 0;
      verilogPut_KeyCollapse_3_680 <= 0;
      verilogPut_Data_3_681 <= 0;
      verilogPut_Found_682 <= 0;
      verilogPut_Key_683 <= 0;
      verilogPut_FoundKey_684 <= 0;
      verilogPut_Data_685 <= 0;
      verilogPut_BtreeIndex_686 <= 0;
      verilogPut_StuckIndex_687 <= 0;
      verilogPut_MergeSuccess_688 <= 0;
      verilogPut_index_689 <= 0;
      verilogPut_size_690 <= 0;
      verilogPut_isLeaf_691 <= 0;
      verilogPut_nextFree_692 <= 0;
      verilogPut_Key_0_693 <= 0;
      verilogPut_KeyCompares_0_694 <= 0;
      verilogPut_KeyCollapse_0_695 <= 0;
      verilogPut_Data_0_696 <= 0;
      verilogPut_Key_1_697 <= 0;
      verilogPut_KeyCompares_1_698 <= 0;
      verilogPut_KeyCollapse_1_699 <= 0;
      verilogPut_Data_1_700 <= 0;
      verilogPut_Key_2_701 <= 0;
      verilogPut_KeyCompares_2_702 <= 0;
      verilogPut_KeyCollapse_2_703 <= 0;
      verilogPut_Data_2_704 <= 0;
      verilogPut_Key_3_705 <= 0;
      verilogPut_KeyCompares_3_706 <= 0;
      verilogPut_KeyCollapse_3_707 <= 0;
      verilogPut_Data_3_708 <= 0;
      verilogPut_Found_709 <= 0;
      verilogPut_Key_710 <= 0;
      verilogPut_FoundKey_711 <= 0;
      verilogPut_Data_712 <= 0;
      verilogPut_BtreeIndex_713 <= 0;
      verilogPut_StuckIndex_714 <= 0;
      verilogPut_MergeSuccess_715 <= 0;
      verilogPut_index_716 <= 0;
      verilogPut_size_717 <= 0;
      verilogPut_isLeaf_718 <= 0;
      verilogPut_nextFree_719 <= 0;
      verilogPut_Key_0_720 <= 0;
      verilogPut_KeyCompares_0_721 <= 0;
      verilogPut_KeyCollapse_0_722 <= 0;
      verilogPut_Data_0_723 <= 0;
      verilogPut_Key_1_724 <= 0;
      verilogPut_KeyCompares_1_725 <= 0;
      verilogPut_KeyCollapse_1_726 <= 0;
      verilogPut_Data_1_727 <= 0;
      verilogPut_Key_2_728 <= 0;
      verilogPut_KeyCompares_2_729 <= 0;
      verilogPut_KeyCollapse_2_730 <= 0;
      verilogPut_Data_2_731 <= 0;
      verilogPut_Key_3_732 <= 0;
      verilogPut_KeyCompares_3_733 <= 0;
      verilogPut_KeyCollapse_3_734 <= 0;
      verilogPut_Data_3_735 <= 0;
      verilogPut_Found_736 <= 0;
      verilogPut_Key_737 <= 0;
      verilogPut_FoundKey_738 <= 0;
      verilogPut_Data_739 <= 0;
      verilogPut_BtreeIndex_740 <= 0;
      verilogPut_StuckIndex_741 <= 0;
      verilogPut_MergeSuccess_742 <= 0;
      verilogPut_childKey_743 <= 0;
      verilogPut_childData_744 <= 0;
      verilogPut_indexLeft_745 <= 0;
      verilogPut_indexRight_746 <= 0;
      verilogPut_midKey_747 <= 0;
      verilogPut_root_748 <= 0;
      verilogPut_next_749 <= 0;
      verilogPut_isLeaf_750 <= 0;
      verilogPut_isFree_751 <= 0;
      verilogPut_index_752 <= 0;
      verilogPut_size_753 <= 0;
      verilogPut_isLeaf_754 <= 0;
      verilogPut_nextFree_755 <= 0;
      verilogPut_Key_0_756 <= 0;
      verilogPut_KeyCompares_0_757 <= 0;
      verilogPut_KeyCollapse_0_758 <= 0;
      verilogPut_Data_0_759 <= 0;
      verilogPut_Key_1_760 <= 0;
      verilogPut_KeyCompares_1_761 <= 0;
      verilogPut_KeyCollapse_1_762 <= 0;
      verilogPut_Data_1_763 <= 0;
      verilogPut_Key_2_764 <= 0;
      verilogPut_KeyCompares_2_765 <= 0;
      verilogPut_KeyCollapse_2_766 <= 0;
      verilogPut_Data_2_767 <= 0;
      verilogPut_Key_3_768 <= 0;
      verilogPut_KeyCompares_3_769 <= 0;
      verilogPut_KeyCollapse_3_770 <= 0;
      verilogPut_Data_3_771 <= 0;
      verilogPut_Found_772 <= 0;
      verilogPut_Key_773 <= 0;
      verilogPut_FoundKey_774 <= 0;
      verilogPut_Data_775 <= 0;
      verilogPut_BtreeIndex_776 <= 0;
      verilogPut_StuckIndex_777 <= 0;
      verilogPut_MergeSuccess_778 <= 0;
      verilogPut_position_779 <= 0;
      verilogPut_index_780 <= 0;
      verilogPut_within_781 <= 0;
      verilogPut_isLeaf_782 <= 0;
      verilogPut_index_783 <= 0;
      verilogPut_size_784 <= 0;
      verilogPut_isLeaf_785 <= 0;
      verilogPut_nextFree_786 <= 0;
      verilogPut_Key_0_787 <= 0;
      verilogPut_KeyCompares_0_788 <= 0;
      verilogPut_KeyCollapse_0_789 <= 0;
      verilogPut_Data_0_790 <= 0;
      verilogPut_Key_1_791 <= 0;
      verilogPut_KeyCompares_1_792 <= 0;
      verilogPut_KeyCollapse_1_793 <= 0;
      verilogPut_Data_1_794 <= 0;
      verilogPut_Key_2_795 <= 0;
      verilogPut_KeyCompares_2_796 <= 0;
      verilogPut_KeyCollapse_2_797 <= 0;
      verilogPut_Data_2_798 <= 0;
      verilogPut_Key_3_799 <= 0;
      verilogPut_KeyCompares_3_800 <= 0;
      verilogPut_KeyCollapse_3_801 <= 0;
      verilogPut_Data_3_802 <= 0;
      verilogPut_Found_803 <= 0;
      verilogPut_Key_804 <= 0;
      verilogPut_FoundKey_805 <= 0;
      verilogPut_Data_806 <= 0;
      verilogPut_BtreeIndex_807 <= 0;
      verilogPut_StuckIndex_808 <= 0;
      verilogPut_MergeSuccess_809 <= 0;
      verilogPut_index_810 <= 0;
      verilogPut_size_811 <= 0;
      verilogPut_isLeaf_812 <= 0;
      verilogPut_nextFree_813 <= 0;
      verilogPut_Key_0_814 <= 0;
      verilogPut_KeyCompares_0_815 <= 0;
      verilogPut_KeyCollapse_0_816 <= 0;
      verilogPut_Data_0_817 <= 0;
      verilogPut_Key_1_818 <= 0;
      verilogPut_KeyCompares_1_819 <= 0;
      verilogPut_KeyCollapse_1_820 <= 0;
      verilogPut_Data_1_821 <= 0;
      verilogPut_Key_2_822 <= 0;
      verilogPut_KeyCompares_2_823 <= 0;
      verilogPut_KeyCollapse_2_824 <= 0;
      verilogPut_Data_2_825 <= 0;
      verilogPut_Key_3_826 <= 0;
      verilogPut_KeyCompares_3_827 <= 0;
      verilogPut_KeyCollapse_3_828 <= 0;
      verilogPut_Data_3_829 <= 0;
      verilogPut_Found_830 <= 0;
      verilogPut_Key_831 <= 0;
      verilogPut_FoundKey_832 <= 0;
      verilogPut_Data_833 <= 0;
      verilogPut_BtreeIndex_834 <= 0;
      verilogPut_StuckIndex_835 <= 0;
      verilogPut_MergeSuccess_836 <= 0;
      verilogPut_index_837 <= 0;
      verilogPut_size_838 <= 0;
      verilogPut_isLeaf_839 <= 0;
      verilogPut_nextFree_840 <= 0;
      verilogPut_Key_0_841 <= 0;
      verilogPut_KeyCompares_0_842 <= 0;
      verilogPut_KeyCollapse_0_843 <= 0;
      verilogPut_Data_0_844 <= 0;
      verilogPut_Key_1_845 <= 0;
      verilogPut_KeyCompares_1_846 <= 0;
      verilogPut_KeyCollapse_1_847 <= 0;
      verilogPut_Data_1_848 <= 0;
      verilogPut_Key_2_849 <= 0;
      verilogPut_KeyCompares_2_850 <= 0;
      verilogPut_KeyCollapse_2_851 <= 0;
      verilogPut_Data_2_852 <= 0;
      verilogPut_Key_3_853 <= 0;
      verilogPut_KeyCompares_3_854 <= 0;
      verilogPut_KeyCollapse_3_855 <= 0;
      verilogPut_Data_3_856 <= 0;
      verilogPut_Found_857 <= 0;
      verilogPut_Key_858 <= 0;
      verilogPut_FoundKey_859 <= 0;
      verilogPut_Data_860 <= 0;
      verilogPut_BtreeIndex_861 <= 0;
      verilogPut_StuckIndex_862 <= 0;
      verilogPut_MergeSuccess_863 <= 0;
      verilogPut_childKey_864 <= 0;
      verilogPut_childData_865 <= 0;
      verilogPut_indexLeft_866 <= 0;
      verilogPut_indexRight_867 <= 0;
      verilogPut_midKey_868 <= 0;
      verilogPut_success_869 <= 0;
      verilogPut_test_870 <= 0;
      verilogPut_next_871 <= 0;
      verilogPut_root_872 <= 0;
      verilogPut_isFree_873 <= 0;
      verilogPut_next_874 <= 0;
      verilogPut_root_875 <= 0;
      verilogPut_isFree_876 <= 0;
      verilogPut_index_877 <= 0;
      verilogPut_size_878 <= 0;
      verilogPut_isLeaf_879 <= 0;
      verilogPut_nextFree_880 <= 0;
      verilogPut_Key_0_881 <= 0;
      verilogPut_KeyCompares_0_882 <= 0;
      verilogPut_KeyCollapse_0_883 <= 0;
      verilogPut_Data_0_884 <= 0;
      verilogPut_Key_1_885 <= 0;
      verilogPut_KeyCompares_1_886 <= 0;
      verilogPut_KeyCollapse_1_887 <= 0;
      verilogPut_Data_1_888 <= 0;
      verilogPut_Key_2_889 <= 0;
      verilogPut_KeyCompares_2_890 <= 0;
      verilogPut_KeyCollapse_2_891 <= 0;
      verilogPut_Data_2_892 <= 0;
      verilogPut_Key_3_893 <= 0;
      verilogPut_KeyCompares_3_894 <= 0;
      verilogPut_KeyCollapse_3_895 <= 0;
      verilogPut_Data_3_896 <= 0;
      verilogPut_Found_897 <= 0;
      verilogPut_Key_898 <= 0;
      verilogPut_FoundKey_899 <= 0;
      verilogPut_Data_900 <= 0;
      verilogPut_BtreeIndex_901 <= 0;
      verilogPut_StuckIndex_902 <= 0;
      verilogPut_MergeSuccess_903 <= 0;
      verilogPut_index_904 <= 0;
      verilogPut_size_905 <= 0;
      verilogPut_isLeaf_906 <= 0;
      verilogPut_nextFree_907 <= 0;
      verilogPut_Key_0_908 <= 0;
      verilogPut_KeyCompares_0_909 <= 0;
      verilogPut_KeyCollapse_0_910 <= 0;
      verilogPut_Data_0_911 <= 0;
      verilogPut_Key_1_912 <= 0;
      verilogPut_KeyCompares_1_913 <= 0;
      verilogPut_KeyCollapse_1_914 <= 0;
      verilogPut_Data_1_915 <= 0;
      verilogPut_Key_2_916 <= 0;
      verilogPut_KeyCompares_2_917 <= 0;
      verilogPut_KeyCollapse_2_918 <= 0;
      verilogPut_Data_2_919 <= 0;
      verilogPut_Key_3_920 <= 0;
      verilogPut_KeyCompares_3_921 <= 0;
      verilogPut_KeyCollapse_3_922 <= 0;
      verilogPut_Data_3_923 <= 0;
      verilogPut_Found_924 <= 0;
      verilogPut_Key_925 <= 0;
      verilogPut_FoundKey_926 <= 0;
      verilogPut_Data_927 <= 0;
      verilogPut_BtreeIndex_928 <= 0;
      verilogPut_StuckIndex_929 <= 0;
      verilogPut_MergeSuccess_930 <= 0;
      verilogPut_index_931 <= 0;
      verilogPut_size_932 <= 0;
      verilogPut_isLeaf_933 <= 0;
      verilogPut_nextFree_934 <= 0;
      verilogPut_Key_0_935 <= 0;
      verilogPut_KeyCompares_0_936 <= 0;
      verilogPut_KeyCollapse_0_937 <= 0;
      verilogPut_Data_0_938 <= 0;
      verilogPut_Key_1_939 <= 0;
      verilogPut_KeyCompares_1_940 <= 0;
      verilogPut_KeyCollapse_1_941 <= 0;
      verilogPut_Data_1_942 <= 0;
      verilogPut_Key_2_943 <= 0;
      verilogPut_KeyCompares_2_944 <= 0;
      verilogPut_KeyCollapse_2_945 <= 0;
      verilogPut_Data_2_946 <= 0;
      verilogPut_Key_3_947 <= 0;
      verilogPut_KeyCompares_3_948 <= 0;
      verilogPut_KeyCollapse_3_949 <= 0;
      verilogPut_Data_3_950 <= 0;
      verilogPut_Found_951 <= 0;
      verilogPut_Key_952 <= 0;
      verilogPut_FoundKey_953 <= 0;
      verilogPut_Data_954 <= 0;
      verilogPut_BtreeIndex_955 <= 0;
      verilogPut_StuckIndex_956 <= 0;
      verilogPut_MergeSuccess_957 <= 0;
      verilogPut_childKey_958 <= 0;
      verilogPut_leftChild_959 <= 0;
      verilogPut_rightChild_960 <= 0;
      verilogPut_childData_961 <= 0;
      verilogPut_indexLeft_962 <= 0;
      verilogPut_indexRight_963 <= 0;
      verilogPut_midKey_964 <= 0;
      verilogPut_success_965 <= 0;
      verilogPut_test_966 <= 0;
      verilogPut_next_967 <= 0;
      verilogPut_root_968 <= 0;
      verilogPut_isFree_969 <= 0;
      verilogPut_next_970 <= 0;
      verilogPut_root_971 <= 0;
      verilogPut_isFree_972 <= 0;
      verilogPut_index_973 <= 0;
      verilogPut_size_974 <= 0;
      verilogPut_isLeaf_975 <= 0;
      verilogPut_nextFree_976 <= 0;
      verilogPut_Key_0_977 <= 0;
      verilogPut_KeyCompares_0_978 <= 0;
      verilogPut_KeyCollapse_0_979 <= 0;
      verilogPut_Data_0_980 <= 0;
      verilogPut_Key_1_981 <= 0;
      verilogPut_KeyCompares_1_982 <= 0;
      verilogPut_KeyCollapse_1_983 <= 0;
      verilogPut_Data_1_984 <= 0;
      verilogPut_Key_2_985 <= 0;
      verilogPut_KeyCompares_2_986 <= 0;
      verilogPut_KeyCollapse_2_987 <= 0;
      verilogPut_Data_2_988 <= 0;
      verilogPut_Key_3_989 <= 0;
      verilogPut_KeyCompares_3_990 <= 0;
      verilogPut_KeyCollapse_3_991 <= 0;
      verilogPut_Data_3_992 <= 0;
      verilogPut_Found_993 <= 0;
      verilogPut_Key_994 <= 0;
      verilogPut_FoundKey_995 <= 0;
      verilogPut_Data_996 <= 0;
      verilogPut_BtreeIndex_997 <= 0;
      verilogPut_StuckIndex_998 <= 0;
      verilogPut_MergeSuccess_999 <= 0;
      verilogPut_index_1000 <= 0;
      verilogPut_size_1001 <= 0;
      verilogPut_isLeaf_1002 <= 0;
      verilogPut_nextFree_1003 <= 0;
      verilogPut_Key_0_1004 <= 0;
      verilogPut_KeyCompares_0_1005 <= 0;
      verilogPut_KeyCollapse_0_1006 <= 0;
      verilogPut_Data_0_1007 <= 0;
      verilogPut_Key_1_1008 <= 0;
      verilogPut_KeyCompares_1_1009 <= 0;
      verilogPut_KeyCollapse_1_1010 <= 0;
      verilogPut_Data_1_1011 <= 0;
      verilogPut_Key_2_1012 <= 0;
      verilogPut_KeyCompares_2_1013 <= 0;
      verilogPut_KeyCollapse_2_1014 <= 0;
      verilogPut_Data_2_1015 <= 0;
      verilogPut_Key_3_1016 <= 0;
      verilogPut_KeyCompares_3_1017 <= 0;
      verilogPut_KeyCollapse_3_1018 <= 0;
      verilogPut_Data_3_1019 <= 0;
      verilogPut_Found_1020 <= 0;
      verilogPut_Key_1021 <= 0;
      verilogPut_FoundKey_1022 <= 0;
      verilogPut_Data_1023 <= 0;
      verilogPut_BtreeIndex_1024 <= 0;
      verilogPut_StuckIndex_1025 <= 0;
      verilogPut_MergeSuccess_1026 <= 0;
      verilogPut_childKey_1027 <= 0;
      verilogPut_size_1028 <= 0;
      verilogPut_childData_1029 <= 0;
      verilogPut_indexLeft_1030 <= 0;
      verilogPut_indexRight_1031 <= 0;
      verilogPut_midKey_1032 <= 0;
      verilogPut_success_1033 <= 0;
      verilogPut_test_1034 <= 0;
      verilogPut_next_1035 <= 0;
      verilogPut_root_1036 <= 0;
      verilogPut_isFree_1037 <= 0;
      verilogPut_index_1038 <= 0;
      verilogPut_size_1039 <= 0;
      verilogPut_isLeaf_1040 <= 0;
      verilogPut_nextFree_1041 <= 0;
      verilogPut_Key_0_1042 <= 0;
      verilogPut_KeyCompares_0_1043 <= 0;
      verilogPut_KeyCollapse_0_1044 <= 0;
      verilogPut_Data_0_1045 <= 0;
      verilogPut_Key_1_1046 <= 0;
      verilogPut_KeyCompares_1_1047 <= 0;
      verilogPut_KeyCollapse_1_1048 <= 0;
      verilogPut_Data_1_1049 <= 0;
      verilogPut_Key_2_1050 <= 0;
      verilogPut_KeyCompares_2_1051 <= 0;
      verilogPut_KeyCollapse_2_1052 <= 0;
      verilogPut_Data_2_1053 <= 0;
      verilogPut_Key_3_1054 <= 0;
      verilogPut_KeyCompares_3_1055 <= 0;
      verilogPut_KeyCollapse_3_1056 <= 0;
      verilogPut_Data_3_1057 <= 0;
      verilogPut_Found_1058 <= 0;
      verilogPut_Key_1059 <= 0;
      verilogPut_FoundKey_1060 <= 0;
      verilogPut_Data_1061 <= 0;
      verilogPut_BtreeIndex_1062 <= 0;
      verilogPut_StuckIndex_1063 <= 0;
      verilogPut_MergeSuccess_1064 <= 0;
      verilogPut_index_1065 <= 0;
      verilogPut_size_1066 <= 0;
      verilogPut_isLeaf_1067 <= 0;
      verilogPut_nextFree_1068 <= 0;
      verilogPut_Key_0_1069 <= 0;
      verilogPut_KeyCompares_0_1070 <= 0;
      verilogPut_KeyCollapse_0_1071 <= 0;
      verilogPut_Data_0_1072 <= 0;
      verilogPut_Key_1_1073 <= 0;
      verilogPut_KeyCompares_1_1074 <= 0;
      verilogPut_KeyCollapse_1_1075 <= 0;
      verilogPut_Data_1_1076 <= 0;
      verilogPut_Key_2_1077 <= 0;
      verilogPut_KeyCompares_2_1078 <= 0;
      verilogPut_KeyCollapse_2_1079 <= 0;
      verilogPut_Data_2_1080 <= 0;
      verilogPut_Key_3_1081 <= 0;
      verilogPut_KeyCompares_3_1082 <= 0;
      verilogPut_KeyCollapse_3_1083 <= 0;
      verilogPut_Data_3_1084 <= 0;
      verilogPut_Found_1085 <= 0;
      verilogPut_Key_1086 <= 0;
      verilogPut_FoundKey_1087 <= 0;
      verilogPut_Data_1088 <= 0;
      verilogPut_BtreeIndex_1089 <= 0;
      verilogPut_StuckIndex_1090 <= 0;
      verilogPut_MergeSuccess_1091 <= 0;
      verilogPut_childKey_1092 <= 0;
      verilogPut_size_1093 <= 0;
      verilogPut_childData_1094 <= 0;
      verilogPut_indexLeft_1095 <= 0;
      verilogPut_indexRight_1096 <= 0;
      verilogPut_midKey_1097 <= 0;
      verilogPut_success_1098 <= 0;
      verilogPut_test_1099 <= 0;
      verilogPut_next_1100 <= 0;
      verilogPut_root_1101 <= 0;
      verilogPut_isFree_1102 <= 0;
      verilogPut_index_1103 <= 0;
      verilogPut_size_1104 <= 0;
      verilogPut_isLeaf_1105 <= 0;
      verilogPut_nextFree_1106 <= 0;
      verilogPut_Key_0_1107 <= 0;
      verilogPut_KeyCompares_0_1108 <= 0;
      verilogPut_KeyCollapse_0_1109 <= 0;
      verilogPut_Data_0_1110 <= 0;
      verilogPut_Key_1_1111 <= 0;
      verilogPut_KeyCompares_1_1112 <= 0;
      verilogPut_KeyCollapse_1_1113 <= 0;
      verilogPut_Data_1_1114 <= 0;
      verilogPut_Key_2_1115 <= 0;
      verilogPut_KeyCompares_2_1116 <= 0;
      verilogPut_KeyCollapse_2_1117 <= 0;
      verilogPut_Data_2_1118 <= 0;
      verilogPut_Key_3_1119 <= 0;
      verilogPut_KeyCompares_3_1120 <= 0;
      verilogPut_KeyCollapse_3_1121 <= 0;
      verilogPut_Data_3_1122 <= 0;
      verilogPut_Found_1123 <= 0;
      verilogPut_Key_1124 <= 0;
      verilogPut_FoundKey_1125 <= 0;
      verilogPut_Data_1126 <= 0;
      verilogPut_BtreeIndex_1127 <= 0;
      verilogPut_StuckIndex_1128 <= 0;
      verilogPut_MergeSuccess_1129 <= 0;
      verilogPut_index_1130 <= 0;
      verilogPut_size_1131 <= 0;
      verilogPut_isLeaf_1132 <= 0;
      verilogPut_nextFree_1133 <= 0;
      verilogPut_Key_0_1134 <= 0;
      verilogPut_KeyCompares_0_1135 <= 0;
      verilogPut_KeyCollapse_0_1136 <= 0;
      verilogPut_Data_0_1137 <= 0;
      verilogPut_Key_1_1138 <= 0;
      verilogPut_KeyCompares_1_1139 <= 0;
      verilogPut_KeyCollapse_1_1140 <= 0;
      verilogPut_Data_1_1141 <= 0;
      verilogPut_Key_2_1142 <= 0;
      verilogPut_KeyCompares_2_1143 <= 0;
      verilogPut_KeyCollapse_2_1144 <= 0;
      verilogPut_Data_2_1145 <= 0;
      verilogPut_Key_3_1146 <= 0;
      verilogPut_KeyCompares_3_1147 <= 0;
      verilogPut_KeyCollapse_3_1148 <= 0;
      verilogPut_Data_3_1149 <= 0;
      verilogPut_Found_1150 <= 0;
      verilogPut_Key_1151 <= 0;
      verilogPut_FoundKey_1152 <= 0;
      verilogPut_Data_1153 <= 0;
      verilogPut_BtreeIndex_1154 <= 0;
      verilogPut_StuckIndex_1155 <= 0;
      verilogPut_MergeSuccess_1156 <= 0;
      verilogPut_childKey_1157 <= 0;
      verilogPut_childData_1158 <= 0;
      verilogPut_indexLeft_1159 <= 0;
      verilogPut_indexRight_1160 <= 0;
      verilogPut_midKey_1161 <= 0;
      verilogPut_success_1162 <= 0;
      verilogPut_test_1163 <= 0;
      verilogPut_next_1164 <= 0;
      verilogPut_root_1165 <= 0;
      verilogPut_isFree_1166 <= 0;
      verilogPut_index_1167 <= 0;
      verilogPut_size_1168 <= 0;
      verilogPut_isLeaf_1169 <= 0;
      verilogPut_nextFree_1170 <= 0;
      verilogPut_Key_0_1171 <= 0;
      verilogPut_KeyCompares_0_1172 <= 0;
      verilogPut_KeyCollapse_0_1173 <= 0;
      verilogPut_Data_0_1174 <= 0;
      verilogPut_Key_1_1175 <= 0;
      verilogPut_KeyCompares_1_1176 <= 0;
      verilogPut_KeyCollapse_1_1177 <= 0;
      verilogPut_Data_1_1178 <= 0;
      verilogPut_Key_2_1179 <= 0;
      verilogPut_KeyCompares_2_1180 <= 0;
      verilogPut_KeyCollapse_2_1181 <= 0;
      verilogPut_Data_2_1182 <= 0;
      verilogPut_Key_3_1183 <= 0;
      verilogPut_KeyCompares_3_1184 <= 0;
      verilogPut_KeyCollapse_3_1185 <= 0;
      verilogPut_Data_3_1186 <= 0;
      verilogPut_Found_1187 <= 0;
      verilogPut_Key_1188 <= 0;
      verilogPut_FoundKey_1189 <= 0;
      verilogPut_Data_1190 <= 0;
      verilogPut_BtreeIndex_1191 <= 0;
      verilogPut_StuckIndex_1192 <= 0;
      verilogPut_MergeSuccess_1193 <= 0;
      verilogPut_index_1194 <= 0;
      verilogPut_size_1195 <= 0;
      verilogPut_isLeaf_1196 <= 0;
      verilogPut_nextFree_1197 <= 0;
      verilogPut_Key_0_1198 <= 0;
      verilogPut_KeyCompares_0_1199 <= 0;
      verilogPut_KeyCollapse_0_1200 <= 0;
      verilogPut_Data_0_1201 <= 0;
      verilogPut_Key_1_1202 <= 0;
      verilogPut_KeyCompares_1_1203 <= 0;
      verilogPut_KeyCollapse_1_1204 <= 0;
      verilogPut_Data_1_1205 <= 0;
      verilogPut_Key_2_1206 <= 0;
      verilogPut_KeyCompares_2_1207 <= 0;
      verilogPut_KeyCollapse_2_1208 <= 0;
      verilogPut_Data_2_1209 <= 0;
      verilogPut_Key_3_1210 <= 0;
      verilogPut_KeyCompares_3_1211 <= 0;
      verilogPut_KeyCollapse_3_1212 <= 0;
      verilogPut_Data_3_1213 <= 0;
      verilogPut_Found_1214 <= 0;
      verilogPut_Key_1215 <= 0;
      verilogPut_FoundKey_1216 <= 0;
      verilogPut_Data_1217 <= 0;
      verilogPut_BtreeIndex_1218 <= 0;
      verilogPut_StuckIndex_1219 <= 0;
      verilogPut_MergeSuccess_1220 <= 0;
      verilogPut_childKey_1221 <= 0;
      verilogPut_leftChild_1222 <= 0;
      verilogPut_rightChild_1223 <= 0;
      verilogPut_childData_1224 <= 0;
      verilogPut_indexLeft_1225 <= 0;
      verilogPut_indexRight_1226 <= 0;
      verilogPut_midKey_1227 <= 0;
      verilogPut_success_1228 <= 0;
      verilogPut_test_1229 <= 0;
      verilogPut_next_1230 <= 0;
      verilogPut_root_1231 <= 0;
      verilogPut_isFree_1232 <= 0;
      verilogPut_index_1233 <= 0;
      verilogPut_size_1234 <= 0;
      verilogPut_isLeaf_1235 <= 0;
      verilogPut_nextFree_1236 <= 0;
      verilogPut_Key_0_1237 <= 0;
      verilogPut_KeyCompares_0_1238 <= 0;
      verilogPut_KeyCollapse_0_1239 <= 0;
      verilogPut_Data_0_1240 <= 0;
      verilogPut_Key_1_1241 <= 0;
      verilogPut_KeyCompares_1_1242 <= 0;
      verilogPut_KeyCollapse_1_1243 <= 0;
      verilogPut_Data_1_1244 <= 0;
      verilogPut_Key_2_1245 <= 0;
      verilogPut_KeyCompares_2_1246 <= 0;
      verilogPut_KeyCollapse_2_1247 <= 0;
      verilogPut_Data_2_1248 <= 0;
      verilogPut_Key_3_1249 <= 0;
      verilogPut_KeyCompares_3_1250 <= 0;
      verilogPut_KeyCollapse_3_1251 <= 0;
      verilogPut_Data_3_1252 <= 0;
      verilogPut_Found_1253 <= 0;
      verilogPut_Key_1254 <= 0;
      verilogPut_FoundKey_1255 <= 0;
      verilogPut_Data_1256 <= 0;
      verilogPut_BtreeIndex_1257 <= 0;
      verilogPut_StuckIndex_1258 <= 0;
      verilogPut_MergeSuccess_1259 <= 0;
      verilogPut_index_1260 <= 0;
      verilogPut_size_1261 <= 0;
      verilogPut_isLeaf_1262 <= 0;
      verilogPut_nextFree_1263 <= 0;
      verilogPut_Key_0_1264 <= 0;
      verilogPut_KeyCompares_0_1265 <= 0;
      verilogPut_KeyCollapse_0_1266 <= 0;
      verilogPut_Data_0_1267 <= 0;
      verilogPut_Key_1_1268 <= 0;
      verilogPut_KeyCompares_1_1269 <= 0;
      verilogPut_KeyCollapse_1_1270 <= 0;
      verilogPut_Data_1_1271 <= 0;
      verilogPut_Key_2_1272 <= 0;
      verilogPut_KeyCompares_2_1273 <= 0;
      verilogPut_KeyCollapse_2_1274 <= 0;
      verilogPut_Data_2_1275 <= 0;
      verilogPut_Key_3_1276 <= 0;
      verilogPut_KeyCompares_3_1277 <= 0;
      verilogPut_KeyCollapse_3_1278 <= 0;
      verilogPut_Data_3_1279 <= 0;
      verilogPut_Found_1280 <= 0;
      verilogPut_Key_1281 <= 0;
      verilogPut_FoundKey_1282 <= 0;
      verilogPut_Data_1283 <= 0;
      verilogPut_BtreeIndex_1284 <= 0;
      verilogPut_StuckIndex_1285 <= 0;
      verilogPut_MergeSuccess_1286 <= 0;
      verilogPut_childKey_1287 <= 0;
      verilogPut_childData_1288 <= 0;
      verilogPut_indexLeft_1289 <= 0;
      verilogPut_indexRight_1290 <= 0;
      verilogPut_midKey_1291 <= 0;
      verilogPut_success_1292 <= 0;
      verilogPut_test_1293 <= 0;
      verilogPut_next_1294 <= 0;
      verilogPut_root_1295 <= 0;
      verilogPut_isFree_1296 <= 0;
      verilogPut_index_1297 <= 0;
      verilogPut_size_1298 <= 0;
      verilogPut_isLeaf_1299 <= 0;
      verilogPut_nextFree_1300 <= 0;
      verilogPut_Key_0_1301 <= 0;
      verilogPut_KeyCompares_0_1302 <= 0;
      verilogPut_KeyCollapse_0_1303 <= 0;
      verilogPut_Data_0_1304 <= 0;
      verilogPut_Key_1_1305 <= 0;
      verilogPut_KeyCompares_1_1306 <= 0;
      verilogPut_KeyCollapse_1_1307 <= 0;
      verilogPut_Data_1_1308 <= 0;
      verilogPut_Key_2_1309 <= 0;
      verilogPut_KeyCompares_2_1310 <= 0;
      verilogPut_KeyCollapse_2_1311 <= 0;
      verilogPut_Data_2_1312 <= 0;
      verilogPut_Key_3_1313 <= 0;
      verilogPut_KeyCompares_3_1314 <= 0;
      verilogPut_KeyCollapse_3_1315 <= 0;
      verilogPut_Data_3_1316 <= 0;
      verilogPut_Found_1317 <= 0;
      verilogPut_Key_1318 <= 0;
      verilogPut_FoundKey_1319 <= 0;
      verilogPut_Data_1320 <= 0;
      verilogPut_BtreeIndex_1321 <= 0;
      verilogPut_StuckIndex_1322 <= 0;
      verilogPut_MergeSuccess_1323 <= 0;
      verilogPut_index_1324 <= 0;
      verilogPut_size_1325 <= 0;
      verilogPut_isLeaf_1326 <= 0;
      verilogPut_nextFree_1327 <= 0;
      verilogPut_Key_0_1328 <= 0;
      verilogPut_KeyCompares_0_1329 <= 0;
      verilogPut_KeyCollapse_0_1330 <= 0;
      verilogPut_Data_0_1331 <= 0;
      verilogPut_Key_1_1332 <= 0;
      verilogPut_KeyCompares_1_1333 <= 0;
      verilogPut_KeyCollapse_1_1334 <= 0;
      verilogPut_Data_1_1335 <= 0;
      verilogPut_Key_2_1336 <= 0;
      verilogPut_KeyCompares_2_1337 <= 0;
      verilogPut_KeyCollapse_2_1338 <= 0;
      verilogPut_Data_2_1339 <= 0;
      verilogPut_Key_3_1340 <= 0;
      verilogPut_KeyCompares_3_1341 <= 0;
      verilogPut_KeyCollapse_3_1342 <= 0;
      verilogPut_Data_3_1343 <= 0;
      verilogPut_Found_1344 <= 0;
      verilogPut_Key_1345 <= 0;
      verilogPut_FoundKey_1346 <= 0;
      verilogPut_Data_1347 <= 0;
      verilogPut_BtreeIndex_1348 <= 0;
      verilogPut_StuckIndex_1349 <= 0;
      verilogPut_MergeSuccess_1350 <= 0;
      verilogPut_childKey_1351 <= 0;
      verilogPut_leftChild_1352 <= 0;
      verilogPut_rightChild_1353 <= 0;
      verilogPut_childData_1354 <= 0;
      verilogPut_indexLeft_1355 <= 0;
      verilogPut_indexRight_1356 <= 0;
      verilogPut_midKey_1357 <= 0;
      verilogPut_success_1358 <= 0;
      verilogPut_test_1359 <= 0;
      verilogPut_next_1360 <= 0;
      verilogPut_root_1361 <= 0;
      verilogPut_isFree_1362 <= 0;
      verilogPut_index_1363 <= 0;
      verilogPut_size_1364 <= 0;
      verilogPut_isLeaf_1365 <= 0;
      verilogPut_nextFree_1366 <= 0;
      verilogPut_Key_0_1367 <= 0;
      verilogPut_KeyCompares_0_1368 <= 0;
      verilogPut_KeyCollapse_0_1369 <= 0;
      verilogPut_Data_0_1370 <= 0;
      verilogPut_Key_1_1371 <= 0;
      verilogPut_KeyCompares_1_1372 <= 0;
      verilogPut_KeyCollapse_1_1373 <= 0;
      verilogPut_Data_1_1374 <= 0;
      verilogPut_Key_2_1375 <= 0;
      verilogPut_KeyCompares_2_1376 <= 0;
      verilogPut_KeyCollapse_2_1377 <= 0;
      verilogPut_Data_2_1378 <= 0;
      verilogPut_Key_3_1379 <= 0;
      verilogPut_KeyCompares_3_1380 <= 0;
      verilogPut_KeyCollapse_3_1381 <= 0;
      verilogPut_Data_3_1382 <= 0;
      verilogPut_Found_1383 <= 0;
      verilogPut_Key_1384 <= 0;
      verilogPut_FoundKey_1385 <= 0;
      verilogPut_Data_1386 <= 0;
      verilogPut_BtreeIndex_1387 <= 0;
      verilogPut_StuckIndex_1388 <= 0;
      verilogPut_MergeSuccess_1389 <= 0;
      verilogPut_index_1390 <= 0;
      verilogPut_size_1391 <= 0;
      verilogPut_isLeaf_1392 <= 0;
      verilogPut_nextFree_1393 <= 0;
      verilogPut_Key_0_1394 <= 0;
      verilogPut_KeyCompares_0_1395 <= 0;
      verilogPut_KeyCollapse_0_1396 <= 0;
      verilogPut_Data_0_1397 <= 0;
      verilogPut_Key_1_1398 <= 0;
      verilogPut_KeyCompares_1_1399 <= 0;
      verilogPut_KeyCollapse_1_1400 <= 0;
      verilogPut_Data_1_1401 <= 0;
      verilogPut_Key_2_1402 <= 0;
      verilogPut_KeyCompares_2_1403 <= 0;
      verilogPut_KeyCollapse_2_1404 <= 0;
      verilogPut_Data_2_1405 <= 0;
      verilogPut_Key_3_1406 <= 0;
      verilogPut_KeyCompares_3_1407 <= 0;
      verilogPut_KeyCollapse_3_1408 <= 0;
      verilogPut_Data_3_1409 <= 0;
      verilogPut_Found_1410 <= 0;
      verilogPut_Key_1411 <= 0;
      verilogPut_FoundKey_1412 <= 0;
      verilogPut_Data_1413 <= 0;
      verilogPut_BtreeIndex_1414 <= 0;
      verilogPut_StuckIndex_1415 <= 0;
      verilogPut_MergeSuccess_1416 <= 0;
      verilogPut_childKey_1417 <= 0;
      verilogPut_childData_1418 <= 0;
      verilogPut_indexLeft_1419 <= 0;
      verilogPut_indexRight_1420 <= 0;
      verilogPut_midKey_1421 <= 0;
      verilogPut_success_1422 <= 0;
      verilogPut_test_1423 <= 0;
      verilogPut_next_1424 <= 0;
      verilogPut_root_1425 <= 0;
      verilogPut_isFree_1426 <= 0;
      verilogPut_index_1427 <= 0;
      verilogPut_size_1428 <= 0;
      verilogPut_isLeaf_1429 <= 0;
      verilogPut_nextFree_1430 <= 0;
      verilogPut_Key_0_1431 <= 0;
      verilogPut_KeyCompares_0_1432 <= 0;
      verilogPut_KeyCollapse_0_1433 <= 0;
      verilogPut_Data_0_1434 <= 0;
      verilogPut_Key_1_1435 <= 0;
      verilogPut_KeyCompares_1_1436 <= 0;
      verilogPut_KeyCollapse_1_1437 <= 0;
      verilogPut_Data_1_1438 <= 0;
      verilogPut_Key_2_1439 <= 0;
      verilogPut_KeyCompares_2_1440 <= 0;
      verilogPut_KeyCollapse_2_1441 <= 0;
      verilogPut_Data_2_1442 <= 0;
      verilogPut_Key_3_1443 <= 0;
      verilogPut_KeyCompares_3_1444 <= 0;
      verilogPut_KeyCollapse_3_1445 <= 0;
      verilogPut_Data_3_1446 <= 0;
      verilogPut_Found_1447 <= 0;
      verilogPut_Key_1448 <= 0;
      verilogPut_FoundKey_1449 <= 0;
      verilogPut_Data_1450 <= 0;
      verilogPut_BtreeIndex_1451 <= 0;
      verilogPut_StuckIndex_1452 <= 0;
      verilogPut_MergeSuccess_1453 <= 0;
      verilogPut_index_1454 <= 0;
      verilogPut_size_1455 <= 0;
      verilogPut_isLeaf_1456 <= 0;
      verilogPut_nextFree_1457 <= 0;
      verilogPut_Key_0_1458 <= 0;
      verilogPut_KeyCompares_0_1459 <= 0;
      verilogPut_KeyCollapse_0_1460 <= 0;
      verilogPut_Data_0_1461 <= 0;
      verilogPut_Key_1_1462 <= 0;
      verilogPut_KeyCompares_1_1463 <= 0;
      verilogPut_KeyCollapse_1_1464 <= 0;
      verilogPut_Data_1_1465 <= 0;
      verilogPut_Key_2_1466 <= 0;
      verilogPut_KeyCompares_2_1467 <= 0;
      verilogPut_KeyCollapse_2_1468 <= 0;
      verilogPut_Data_2_1469 <= 0;
      verilogPut_Key_3_1470 <= 0;
      verilogPut_KeyCompares_3_1471 <= 0;
      verilogPut_KeyCollapse_3_1472 <= 0;
      verilogPut_Data_3_1473 <= 0;
      verilogPut_Found_1474 <= 0;
      verilogPut_Key_1475 <= 0;
      verilogPut_FoundKey_1476 <= 0;
      verilogPut_Data_1477 <= 0;
      verilogPut_BtreeIndex_1478 <= 0;
      verilogPut_StuckIndex_1479 <= 0;
      verilogPut_MergeSuccess_1480 <= 0;
      verilogPut_childKey_1481 <= 0;
      verilogPut_leftChild_1482 <= 0;
      verilogPut_rightChild_1483 <= 0;
      verilogPut_childData_1484 <= 0;
      verilogPut_indexLeft_1485 <= 0;
      verilogPut_indexRight_1486 <= 0;
      verilogPut_midKey_1487 <= 0;
      verilogPut_success_1488 <= 0;
      verilogPut_test_1489 <= 0;
      verilogPut_next_1490 <= 0;
      verilogPut_root_1491 <= 0;
      verilogPut_isFree_1492 <= 0;
      stuckIsLeaf_19_requestedAt <= -1;
      stuckIsLeaf_20_requestedAt <= -1;
      stuckIsFree_23_requestedAt <= -1;
      freeNext_21_requestedAt <= -1;
      freeNext_22_requestedAt <= -1;
      stuckSize_17_requestedAt <= -1;
      stuckSize_18_requestedAt <= -1;
      stuckKeys_0_1_requestedAt <= -1;
      stuckKeys_0_2_requestedAt <= -1;
      stuckKeys_1_5_requestedAt <= -1;
      stuckKeys_1_6_requestedAt <= -1;
      stuckKeys_2_9_requestedAt <= -1;
      stuckKeys_2_10_requestedAt <= -1;
      stuckKeys_3_13_requestedAt <= -1;
      stuckKeys_3_14_requestedAt <= -1;
      stuckData_0_3_requestedAt <= -1;
      stuckData_0_4_requestedAt <= -1;
      stuckData_1_7_requestedAt <= -1;
      stuckData_1_8_requestedAt <= -1;
      stuckData_2_11_requestedAt <= -1;
      stuckData_2_12_requestedAt <= -1;
      stuckData_3_15_requestedAt <= -1;
      stuckData_3_16_requestedAt <= -1;
    end
    else begin                                   // Run the process in full parallel
      case(verilogPut_pc)
        0: begin
          verilogPut_k_0 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1: begin
          verilogPut_d_1 <= 11;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        2: begin
          verilogPut_BtreeIndex_110 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        3: begin
          verilogPut_index_86 <= verilogPut_BtreeIndex_110;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        4: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_86;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_86;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_86;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_86;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_86;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_86;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_86;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_86;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_86;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_86;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        5: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        6: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        7: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        8: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        9: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        10: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        11: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        12: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        13: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        14: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        15: begin
          verilogPut_size_87 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_88 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_90 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_93 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_94 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_97 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_98 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_101 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_102 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_105 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        16: begin
          if (verilogPut_isLeaf_88 == 0) begin
            verilogPut_pc <= 23;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        17: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 == verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 == verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 == verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 == verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        18: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        19: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        20: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Key_107 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Key_107 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Key_107 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Key_107 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        21: begin
          verilogPut_pc <= 29;
        end
        22: begin
          verilogPut_pc <= 29;
        end
        23: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 <= verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 >  verilogPut_Key_0_90 && verilogPut_k_0 <= verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 >  verilogPut_Key_1_94 && verilogPut_k_0 <= verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 >  verilogPut_Key_2_98 && verilogPut_k_0 <= verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        24: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        25: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        26: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_FoundKey_108 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_FoundKey_108 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_FoundKey_108 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_FoundKey_108 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
            case (verilogPut_size_87)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        27: begin
          verilogPut_BtreeIndex_110 <= verilogPut_Data_109;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        28: begin
          verilogPut_pc <= 3;
        end
        29: begin
          if (verilogPut_Found_106 == 0) begin
            verilogPut_pc <= 32;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        30: begin
          if (verilogPut_StuckIndex_111 == verilogPut_size_87) begin
            verilogPut_size_87 <= verilogPut_size_87+1;
          end
          case (verilogPut_StuckIndex_111)
            0: begin
              verilogPut_Key_0_90 <= verilogPut_k_0;
              verilogPut_Data_0_93 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_94 <= verilogPut_k_0;
              verilogPut_Data_1_97 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_98 <= verilogPut_k_0;
              verilogPut_Data_2_101 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_102 <= verilogPut_k_0;
              verilogPut_Data_3_105 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        31: begin
          verilogPut_pc <= 43;
        end
        32: begin
          verilogPut_notFull_119 <= verilogPut_size_87< 4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        33: begin
          if (verilogPut_notFull_119 == 0) begin
            verilogPut_pc <= 42;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        34: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 <= verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 >  verilogPut_Key_0_90 && verilogPut_k_0 <= verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 >  verilogPut_Key_1_94 && verilogPut_k_0 <= verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 >  verilogPut_Key_2_98 && verilogPut_k_0 <= verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        35: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        36: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        37: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_FoundKey_108 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_FoundKey_108 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_FoundKey_108 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_FoundKey_108 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
            case (verilogPut_size_87)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        38: begin
          verilogPut_size_87 <= verilogPut_size_87+1;
          if (3 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_3_102 <= verilogPut_Key_2_98;
            verilogPut_Data_3_105 <= verilogPut_Data_2_101;
          end
          if (2 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_2_98 <= verilogPut_Key_1_94;
            verilogPut_Data_2_101 <= verilogPut_Data_1_97;
          end
          if (1 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_1_94 <= verilogPut_Key_0_90;
            verilogPut_Data_1_97 <= verilogPut_Data_0_93;
          end
          case (verilogPut_StuckIndex_111)
            0: begin
              verilogPut_Key_0_90 <= verilogPut_k_0;
              verilogPut_Data_0_93 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_94 <= verilogPut_k_0;
              verilogPut_Data_1_97 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_98 <= verilogPut_k_0;
              verilogPut_Data_2_101 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_102 <= verilogPut_k_0;
              verilogPut_Data_3_105 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        39: begin
          verilogPut_Found_106 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        40: begin
          verilogPut_pc <= verilogPut_pc + 1;
        end
        41: begin
          verilogPut_pc <= 43;
        end
        42: begin
          verilogPut_pc <= 53;
        end
        43: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_86;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_87;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_86;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_90;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_86;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_93;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_86;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_94;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_86;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_97;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_86;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_98;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_86;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_101;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_86;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_102;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_86;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_105;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        44: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        45: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        46: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        47: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        48: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        49: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        50: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        51: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        52: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        53: begin
          if (verilogPut_Found_106 >  0) begin
            verilogPut_pc <= 671;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        54: begin
          if (verilogPut_BtreeIndex_110 == 0) begin
            verilogPut_pc <= 56;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        55: begin
          verilogPut_pc <= 185;
        end
        56: begin
          verilogPut_index_120 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        57: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_120;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_120;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_120;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_120;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_120;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_120;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_120;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_120;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_120;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_120;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        58: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        59: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        60: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        61: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        62: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        63: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        64: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        65: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        66: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        67: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        68: begin
          verilogPut_size_121 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_122 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_124 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_127 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_128 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_131 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_132 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_135 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_136 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_139 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        69: begin
          if (verilogPut_size_121 < 4) begin
            verilogPut_pc <= 133;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        70: begin
          verilogPut_Key_0_151 <= verilogPut_Key_0_124;
          verilogPut_Data_0_154 <= verilogPut_Data_0_127;
          verilogPut_Key_1_155 <= verilogPut_Key_1_128;
          verilogPut_Data_1_158 <= verilogPut_Data_1_131;
          verilogPut_size_148 <= 2;
          verilogPut_Key_0_178 <= verilogPut_Key_2_132;
          verilogPut_Data_0_181 <= verilogPut_Data_2_135;
          verilogPut_Key_1_182 <= verilogPut_Key_3_136;
          verilogPut_Data_1_185 <= verilogPut_Data_3_139;
          verilogPut_size_175 <= 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        71: begin
          verilogPut_root_209 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        72: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_209;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        73: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        74: begin
          verilogPut_indexLeft_201 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        75: begin
          if (verilogPut_indexLeft_201 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_211 <= 1;
          verilogPut_isFree_212 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        76: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexLeft_201;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexLeft_201;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_211;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_201;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_212;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        77: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        78: begin
          verilogPut_next_210 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        79: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_209;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_210;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        80: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        81: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        82: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        83: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexLeft_201;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_148;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexLeft_201;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_151;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexLeft_201;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_154;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexLeft_201;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_155;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexLeft_201;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_158;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexLeft_201;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_159;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexLeft_201;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_162;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexLeft_201;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_163;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexLeft_201;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_166;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        84: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        85: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        86: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        87: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        88: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        89: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        90: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        91: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        92: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        93: begin
          verilogPut_root_213 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        94: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_213;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        95: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        96: begin
          verilogPut_indexRight_202 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        97: begin
          if (verilogPut_indexRight_202 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_215 <= 1;
          verilogPut_isFree_216 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        98: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexRight_202;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexRight_202;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_215;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_202;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_216;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        99: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        100: begin
          verilogPut_next_214 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        101: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_213;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_214;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        102: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        103: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        104: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        105: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexRight_202;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_175;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexRight_202;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_178;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexRight_202;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_181;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexRight_202;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_182;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexRight_202;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_185;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexRight_202;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_186;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexRight_202;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_189;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexRight_202;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_190;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexRight_202;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_193;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        106: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        107: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        108: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        109: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        110: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        111: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        112: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        113: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        114: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        115: begin
          case (verilogPut_size_148)
            1: begin
              verilogPut_Key_168 <= verilogPut_Key_0_151;
              verilogPut_Data_170 <= verilogPut_Data_0_154;
            end
            2: begin
              verilogPut_Key_168 <= verilogPut_Key_1_155;
              verilogPut_Data_170 <= verilogPut_Data_1_158;
            end
            3: begin
              verilogPut_Key_168 <= verilogPut_Key_2_159;
              verilogPut_Data_170 <= verilogPut_Data_2_162;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        116: begin
          verilogPut_Key_195 <= verilogPut_Key_0_178;
          verilogPut_Data_197 <= verilogPut_Data_0_181;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        117: begin
          verilogPut_midKey_203 <= (verilogPut_Key_168 + verilogPut_Key_195) / 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        118: begin
          verilogPut_size_121 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        119: begin
          case (verilogPut_size_121)
            0: begin
              verilogPut_Key_0_124 <= verilogPut_midKey_203;
              verilogPut_Data_0_127 <= verilogPut_indexLeft_201;
            end
            1: begin
              verilogPut_Key_1_128 <= verilogPut_midKey_203;
              verilogPut_Data_1_131 <= verilogPut_indexLeft_201;
            end
            2: begin
              verilogPut_Key_2_132 <= verilogPut_midKey_203;
              verilogPut_Data_2_135 <= verilogPut_indexLeft_201;
            end
            3: begin
              verilogPut_Key_3_136 <= verilogPut_midKey_203;
              verilogPut_Data_3_139 <= verilogPut_indexLeft_201;
            end
          endcase
          verilogPut_size_121 <= verilogPut_size_121+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        120: begin
          case (verilogPut_size_121)
            0: begin
              verilogPut_Key_0_124 <= verilogPut_midKey_203;
              verilogPut_Data_0_127 <= verilogPut_indexRight_202;
            end
            1: begin
              verilogPut_Key_1_128 <= verilogPut_midKey_203;
              verilogPut_Data_1_131 <= verilogPut_indexRight_202;
            end
            2: begin
              verilogPut_Key_2_132 <= verilogPut_midKey_203;
              verilogPut_Data_2_135 <= verilogPut_indexRight_202;
            end
            3: begin
              verilogPut_Key_3_136 <= verilogPut_midKey_203;
              verilogPut_Data_3_139 <= verilogPut_indexRight_202;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        121: begin
          verilogPut_isLeaf_122 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        122: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_120;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_121;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_index_120;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_122;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_120;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_124;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_120;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_127;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_120;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_128;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_120;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_131;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_120;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_132;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_120;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_135;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_120;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_136;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_120;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_139;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        123: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        124: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        125: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        126: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        127: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        128: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        129: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        130: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        131: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        132: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        133: begin
          verilogPut_BtreeIndex_110 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        134: begin
          verilogPut_index_86 <= verilogPut_BtreeIndex_110;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        135: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_86;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_86;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_86;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_86;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_86;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_86;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_86;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_86;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_86;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_86;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        136: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        137: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        138: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        139: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        140: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        141: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        142: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        143: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        144: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        145: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        146: begin
          verilogPut_size_87 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_88 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_90 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_93 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_94 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_97 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_98 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_101 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_102 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_105 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        147: begin
          if (verilogPut_isLeaf_88 == 0) begin
            verilogPut_pc <= 154;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        148: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 == verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 == verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 == verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 == verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        149: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        150: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        151: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Key_107 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Key_107 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Key_107 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Key_107 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        152: begin
          verilogPut_pc <= 160;
        end
        153: begin
          verilogPut_pc <= 160;
        end
        154: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 <= verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 >  verilogPut_Key_0_90 && verilogPut_k_0 <= verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 >  verilogPut_Key_1_94 && verilogPut_k_0 <= verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 >  verilogPut_Key_2_98 && verilogPut_k_0 <= verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        155: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        156: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        157: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_FoundKey_108 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_FoundKey_108 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_FoundKey_108 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_FoundKey_108 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
            case (verilogPut_size_87)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        158: begin
          verilogPut_BtreeIndex_110 <= verilogPut_Data_109;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        159: begin
          verilogPut_pc <= 134;
        end
        160: begin
          if (verilogPut_Found_106 == 0) begin
            verilogPut_pc <= 163;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        161: begin
          if (verilogPut_StuckIndex_111 == verilogPut_size_87) begin
            verilogPut_size_87 <= verilogPut_size_87+1;
          end
          case (verilogPut_StuckIndex_111)
            0: begin
              verilogPut_Key_0_90 <= verilogPut_k_0;
              verilogPut_Data_0_93 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_94 <= verilogPut_k_0;
              verilogPut_Data_1_97 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_98 <= verilogPut_k_0;
              verilogPut_Data_2_101 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_102 <= verilogPut_k_0;
              verilogPut_Data_3_105 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        162: begin
          verilogPut_pc <= 174;
        end
        163: begin
          verilogPut_notFull_218 <= verilogPut_size_87< 4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        164: begin
          if (verilogPut_notFull_218 == 0) begin
            verilogPut_pc <= 173;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        165: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 <= verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 >  verilogPut_Key_0_90 && verilogPut_k_0 <= verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 >  verilogPut_Key_1_94 && verilogPut_k_0 <= verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 >  verilogPut_Key_2_98 && verilogPut_k_0 <= verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        166: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        167: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        168: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_FoundKey_108 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_FoundKey_108 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_FoundKey_108 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_FoundKey_108 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
            case (verilogPut_size_87)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        169: begin
          verilogPut_size_87 <= verilogPut_size_87+1;
          if (3 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_3_102 <= verilogPut_Key_2_98;
            verilogPut_Data_3_105 <= verilogPut_Data_2_101;
          end
          if (2 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_2_98 <= verilogPut_Key_1_94;
            verilogPut_Data_2_101 <= verilogPut_Data_1_97;
          end
          if (1 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_1_94 <= verilogPut_Key_0_90;
            verilogPut_Data_1_97 <= verilogPut_Data_0_93;
          end
          case (verilogPut_StuckIndex_111)
            0: begin
              verilogPut_Key_0_90 <= verilogPut_k_0;
              verilogPut_Data_0_93 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_94 <= verilogPut_k_0;
              verilogPut_Data_1_97 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_98 <= verilogPut_k_0;
              verilogPut_Data_2_101 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_102 <= verilogPut_k_0;
              verilogPut_Data_3_105 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        170: begin
          verilogPut_Found_106 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        171: begin
          verilogPut_pc <= verilogPut_pc + 1;
        end
        172: begin
          verilogPut_pc <= 174;
        end
        173: begin
          verilogPut_pc <= 184;
        end
        174: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_86;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_87;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_86;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_90;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_86;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_93;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_86;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_94;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_86;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_97;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_86;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_98;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_86;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_101;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_86;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_102;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_86;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_105;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        175: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        176: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        177: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        178: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        179: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        180: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        181: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        182: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        183: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        184: begin
          verilogPut_pc <= 671;
        end
        185: begin
          verilogPut_index_2 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        186: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_2;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_2;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_2;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_2;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_2;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_2;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_2;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_2;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_2;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_2;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        187: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        188: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        189: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        190: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        191: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        192: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        193: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        194: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        195: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        196: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        197: begin
          verilogPut_size_3 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_4 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_6 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_9 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_16 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_19 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_26 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_29 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_36 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_39 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        198: begin
          verilogPut_full_117 <= verilogPut_size_3>=3 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        199: begin
          if (verilogPut_full_117 == 0) begin
            verilogPut_pc <= 275;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        200: begin
          verilogPut_index_219 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        201: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_219;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_219;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_219;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_219;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_219;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_219;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_219;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_219;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_219;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_219;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        202: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        203: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        204: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        205: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        206: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        207: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        208: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        209: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        210: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        211: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        212: begin
          verilogPut_size_220 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_221 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_223 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_226 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_227 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_230 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_231 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_234 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_235 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_238 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        213: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        214: begin
          verilogPut_Key_0_250 <= verilogPut_Key_0_223;
          verilogPut_Data_0_253 <= verilogPut_Data_0_226;
          verilogPut_size_247 <= 1;
          verilogPut_Data_1_257 <= verilogPut_Data_1_230;
          verilogPut_Key_0_277 <= verilogPut_Key_2_231;
          verilogPut_Data_0_280 <= verilogPut_Data_2_234;
          case (verilogPut_size_220)
            0: begin
              verilogPut_size_274 <= -2;
              verilogPut_Data_1_284 <= verilogPut_Data_3_238;
            end
            1: begin
              verilogPut_size_274 <= -1;
              verilogPut_Data_1_284 <= verilogPut_Data_3_238;
            end
            2: begin
              verilogPut_size_274 <= 0;
              verilogPut_Data_1_284 <= verilogPut_Data_3_238;
            end
            3: begin
              verilogPut_size_274 <= 1;
              verilogPut_Data_1_284 <= verilogPut_Data_3_238;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        215: begin
          verilogPut_root_303 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        216: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_303;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        217: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        218: begin
          verilogPut_indexLeft_300 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        219: begin
          if (verilogPut_indexLeft_300 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_305 <= 0;
          verilogPut_isFree_306 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        220: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexLeft_300;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexLeft_300;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_305;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_300;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_306;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        221: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        222: begin
          verilogPut_next_304 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        223: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_303;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_304;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        224: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        225: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        226: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        227: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexLeft_300;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_247;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexLeft_300;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_250;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexLeft_300;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_253;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexLeft_300;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_254;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexLeft_300;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_257;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexLeft_300;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_258;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexLeft_300;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_261;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexLeft_300;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_262;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexLeft_300;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_265;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        228: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        229: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        230: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        231: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        232: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        233: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        234: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        235: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        236: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        237: begin
          verilogPut_root_307 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        238: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_307;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        239: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        240: begin
          verilogPut_indexRight_301 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        241: begin
          if (verilogPut_indexRight_301 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_309 <= 0;
          verilogPut_isFree_310 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        242: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexRight_301;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexRight_301;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_309;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_301;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_310;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        243: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        244: begin
          verilogPut_next_308 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        245: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_307;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_308;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        246: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        247: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        248: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        249: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexRight_301;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_274;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexRight_301;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_277;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexRight_301;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_280;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexRight_301;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_281;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexRight_301;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_284;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexRight_301;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_285;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexRight_301;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_288;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexRight_301;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_289;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexRight_301;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_292;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        250: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        251: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        252: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        253: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        254: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        255: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        256: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        257: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        258: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        259: begin
          verilogPut_midKey_302 <= verilogPut_Key_1_227;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        260: begin
          verilogPut_size_220 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        261: begin
          case (verilogPut_size_220)
            0: begin
              verilogPut_Key_0_223 <= verilogPut_midKey_302;
              verilogPut_Data_0_226 <= verilogPut_indexLeft_300;
            end
            1: begin
              verilogPut_Key_1_227 <= verilogPut_midKey_302;
              verilogPut_Data_1_230 <= verilogPut_indexLeft_300;
            end
            2: begin
              verilogPut_Key_2_231 <= verilogPut_midKey_302;
              verilogPut_Data_2_234 <= verilogPut_indexLeft_300;
            end
            3: begin
              verilogPut_Key_3_235 <= verilogPut_midKey_302;
              verilogPut_Data_3_238 <= verilogPut_indexLeft_300;
            end
          endcase
          verilogPut_size_220 <= verilogPut_size_220+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        262: begin
          case (verilogPut_size_220)
            0: begin
              verilogPut_Key_0_223 <= verilogPut_midKey_302;
              verilogPut_Data_0_226 <= verilogPut_indexRight_301;
            end
            1: begin
              verilogPut_Key_1_227 <= verilogPut_midKey_302;
              verilogPut_Data_1_230 <= verilogPut_indexRight_301;
            end
            2: begin
              verilogPut_Key_2_231 <= verilogPut_midKey_302;
              verilogPut_Data_2_234 <= verilogPut_indexRight_301;
            end
            3: begin
              verilogPut_Key_3_235 <= verilogPut_midKey_302;
              verilogPut_Data_3_238 <= verilogPut_indexRight_301;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        263: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_219;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_220;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_219;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_223;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_219;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_226;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_219;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_227;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_219;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_230;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_219;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_231;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_219;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_234;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_219;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_235;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_219;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_238;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        264: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        265: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        266: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        267: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        268: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        269: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        270: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        271: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        272: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        273: begin
          verilogPut_pc <= 53;
        end
        274: begin
          verilogPut_pc <= 275;
        end
        275: begin
          verilogPut_parent_114 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        276: begin
          verilogPut_index_2 <= verilogPut_parent_114;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        277: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_2;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_2;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_2;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_2;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_2;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_2;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_2;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_2;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_2;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_2;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        278: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        279: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        280: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        281: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        282: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        283: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        284: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        285: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        286: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        287: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        288: begin
          verilogPut_size_3 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_4 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_6 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_9 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_16 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_19 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_26 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_29 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_36 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_39 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        289: begin
          verilogPut_KeyCompares_0_7 <= verilogPut_k_0 <= verilogPut_Key_0_6 && 0 < verilogPut_size_3;
          verilogPut_KeyCollapse_0_8 <= 0;
          verilogPut_KeyCompares_1_17 <= verilogPut_k_0 >  verilogPut_Key_0_6 && verilogPut_k_0 <= verilogPut_Key_1_16 && 1 < verilogPut_size_3;
          verilogPut_KeyCollapse_1_18 <= 1;
          verilogPut_KeyCompares_2_27 <= verilogPut_k_0 >  verilogPut_Key_1_16 && verilogPut_k_0 <= verilogPut_Key_2_26 && 2 < verilogPut_size_3;
          verilogPut_KeyCollapse_2_28 <= 2;
          verilogPut_KeyCompares_3_37 <= verilogPut_k_0 >  verilogPut_Key_2_26 && verilogPut_k_0 <= verilogPut_Key_3_36 && 3 < verilogPut_size_3;
          verilogPut_KeyCollapse_3_38 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        290: begin
          if (verilogPut_KeyCompares_1_17) begin
            verilogPut_KeyCompares_0_7 <= 1;
            verilogPut_KeyCollapse_0_8 <= verilogPut_KeyCollapse_1_18;
          end
          if (verilogPut_KeyCompares_3_37) begin
            verilogPut_KeyCompares_2_27 <= 1;
            verilogPut_KeyCollapse_2_28 <= verilogPut_KeyCollapse_3_38;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        291: begin
          if (verilogPut_KeyCompares_2_27) begin
            verilogPut_KeyCompares_0_7 <= 1;
            verilogPut_KeyCollapse_0_8 <= verilogPut_KeyCollapse_2_28;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        292: begin
          if (verilogPut_KeyCompares_0_7) begin
            verilogPut_Found_52 <= 1;
            case (verilogPut_KeyCollapse_0_8)
              0: begin
                verilogPut_StuckIndex_57 <= 0;
                verilogPut_FoundKey_54 <= verilogPut_Key_0_6;
                verilogPut_Data_55 <= verilogPut_Data_0_9;
              end
              1: begin
                verilogPut_StuckIndex_57 <= 1;
                verilogPut_FoundKey_54 <= verilogPut_Key_1_16;
                verilogPut_Data_55 <= verilogPut_Data_1_19;
              end
              2: begin
                verilogPut_StuckIndex_57 <= 2;
                verilogPut_FoundKey_54 <= verilogPut_Key_2_26;
                verilogPut_Data_55 <= verilogPut_Data_2_29;
              end
              3: begin
                verilogPut_StuckIndex_57 <= 3;
                verilogPut_FoundKey_54 <= verilogPut_Key_3_36;
                verilogPut_Data_55 <= verilogPut_Data_3_39;
              end
            endcase
          end
          else begin
            verilogPut_Found_52 <= 0;
            case (verilogPut_size_3)
              0: begin
                verilogPut_StuckIndex_57 <= 0;
                verilogPut_Data_55 <= verilogPut_Data_0_9;
              end
              1: begin
                verilogPut_StuckIndex_57 <= 1;
                verilogPut_Data_55 <= verilogPut_Data_1_19;
              end
              2: begin
                verilogPut_StuckIndex_57 <= 2;
                verilogPut_Data_55 <= verilogPut_Data_2_29;
              end
              3: begin
                verilogPut_StuckIndex_57 <= 3;
                verilogPut_Data_55 <= verilogPut_Data_3_39;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        293: begin
          verilogPut_child_113 <= verilogPut_Data_55;
          verilogPut_childInparent_115 <= verilogPut_StuckIndex_57;
          verilogPut_found_116 <= verilogPut_Found_52;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        294: begin
          verilogPut_index_59 <= verilogPut_child_113;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        295: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_59;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_59;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_59;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_59;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_59;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_59;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_59;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_59;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_59;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_59;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        296: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        297: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        298: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        299: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        300: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        301: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        302: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        303: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        304: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        305: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        306: begin
          verilogPut_size_60 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_61 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_63 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_66 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_67 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_70 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_71 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_74 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_75 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_78 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        307: begin
          if (verilogPut_isLeaf_61 == 0) begin
            verilogPut_pc <= 518;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        308: begin
          verilogPut_full_117 <= verilogPut_size_60>=4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        309: begin
          if (verilogPut_full_117 == 0) begin
            verilogPut_pc <= 465;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        310: begin
          if (verilogPut_found_116 == 0) begin
            verilogPut_pc <= 387;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        311: begin
          verilogPut_index_311 <= verilogPut_parent_114;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        312: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_311;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_311;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_311;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_311;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_311;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_311;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_311;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_311;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_311;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_311;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        313: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        314: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        315: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        316: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        317: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        318: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        319: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        320: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        321: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        322: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        323: begin
          verilogPut_size_312 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_313 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_315 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_318 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_319 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_322 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_323 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_326 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_327 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_330 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        324: begin
          case (verilogPut_childInparent_115)
            0: begin
              verilogPut_childKey_419 <= verilogPut_Key_0_315;
              verilogPut_childData_420 <= verilogPut_Data_0_318;
            end
            1: begin
              verilogPut_childKey_419 <= verilogPut_Key_1_319;
              verilogPut_childData_420 <= verilogPut_Data_1_322;
            end
            2: begin
              verilogPut_childKey_419 <= verilogPut_Key_2_323;
              verilogPut_childData_420 <= verilogPut_Data_2_326;
            end
            3: begin
              verilogPut_childKey_419 <= verilogPut_Key_3_327;
              verilogPut_childData_420 <= verilogPut_Data_3_330;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        325: begin
          verilogPut_index_338 <= verilogPut_childData_420;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        326: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_338;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_338;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_338;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_338;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_338;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_338;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_338;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_338;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_338;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_338;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        327: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        328: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        329: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        330: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        331: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        332: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        333: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        334: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        335: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        336: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        337: begin
          verilogPut_size_339 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_340 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_342 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_345 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_346 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_349 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_350 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_353 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_354 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_357 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        338: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        339: begin
          verilogPut_Key_0_369 <= verilogPut_Key_0_342;
          verilogPut_Data_0_372 <= verilogPut_Data_0_345;
          verilogPut_Key_1_373 <= verilogPut_Key_1_346;
          verilogPut_Data_1_376 <= verilogPut_Data_1_349;
          verilogPut_size_366 <= 2;
          verilogPut_Key_0_342 <= verilogPut_Key_2_350;
          verilogPut_Data_0_345 <= verilogPut_Data_2_353;
          verilogPut_Key_1_346 <= verilogPut_Key_3_354;
          verilogPut_Data_1_349 <= verilogPut_Data_3_357;
          verilogPut_size_339 <= 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        340: begin
          verilogPut_root_424 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        341: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_424;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        342: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        343: begin
          verilogPut_indexLeft_421 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        344: begin
          if (verilogPut_indexLeft_421 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_426 <= 1;
          verilogPut_isFree_427 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        345: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexLeft_421;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexLeft_421;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_426;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_421;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_427;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        346: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        347: begin
          verilogPut_next_425 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        348: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_424;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_425;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        349: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        350: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        351: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        352: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_childData_420;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_339;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_childData_420;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_342;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_childData_420;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_345;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_childData_420;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_346;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_childData_420;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_349;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_childData_420;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_350;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_childData_420;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_353;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_childData_420;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_354;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_childData_420;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_357;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        353: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        354: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        355: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        356: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        357: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        358: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        359: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        360: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        361: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        362: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexLeft_421;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_366;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexLeft_421;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_369;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexLeft_421;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_372;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexLeft_421;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_373;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexLeft_421;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_376;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexLeft_421;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_377;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexLeft_421;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_380;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexLeft_421;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_381;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexLeft_421;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_384;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        363: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        364: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        365: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        366: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        367: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        368: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        369: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        370: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        371: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        372: begin
          case (verilogPut_size_366)
            1: begin
              verilogPut_Key_386 <= verilogPut_Key_0_369;
              verilogPut_Data_388 <= verilogPut_Data_0_372;
            end
            2: begin
              verilogPut_Key_386 <= verilogPut_Key_1_373;
              verilogPut_Data_388 <= verilogPut_Data_1_376;
            end
            3: begin
              verilogPut_Key_386 <= verilogPut_Key_2_377;
              verilogPut_Data_388 <= verilogPut_Data_2_380;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        373: begin
          verilogPut_Key_359 <= verilogPut_Key_0_342;
          verilogPut_Data_361 <= verilogPut_Data_0_345;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        374: begin
          verilogPut_midKey_423 <= (verilogPut_Key_386 + verilogPut_Key_359) / 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        375: begin
          verilogPut_size_312 <= verilogPut_size_312+1;
          if (3 > verilogPut_childInparent_115) begin
            verilogPut_Key_3_327 <= verilogPut_Key_2_323;
            verilogPut_Data_3_330 <= verilogPut_Data_2_326;
          end
          if (2 > verilogPut_childInparent_115) begin
            verilogPut_Key_2_323 <= verilogPut_Key_1_319;
            verilogPut_Data_2_326 <= verilogPut_Data_1_322;
          end
          if (1 > verilogPut_childInparent_115) begin
            verilogPut_Key_1_319 <= verilogPut_Key_0_315;
            verilogPut_Data_1_322 <= verilogPut_Data_0_318;
          end
          case (verilogPut_childInparent_115)
            0: begin
              verilogPut_Key_0_315 <= verilogPut_midKey_423;
              verilogPut_Data_0_318 <= verilogPut_indexLeft_421;
            end
            1: begin
              verilogPut_Key_1_319 <= verilogPut_midKey_423;
              verilogPut_Data_1_322 <= verilogPut_indexLeft_421;
            end
            2: begin
              verilogPut_Key_2_323 <= verilogPut_midKey_423;
              verilogPut_Data_2_326 <= verilogPut_indexLeft_421;
            end
            3: begin
              verilogPut_Key_3_327 <= verilogPut_midKey_423;
              verilogPut_Data_3_330 <= verilogPut_indexLeft_421;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        376: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_311;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_312;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_311;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_315;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_311;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_318;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_311;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_319;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_311;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_322;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_311;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_323;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_311;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_326;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_311;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_327;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_311;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_330;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        377: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        378: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        379: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        380: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        381: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        382: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        383: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        384: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        385: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        386: begin
          verilogPut_pc <= 464;
        end
        387: begin
          verilogPut_index_428 <= verilogPut_parent_114;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        388: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_428;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_428;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_428;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_428;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_428;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_428;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_428;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_428;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_428;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_428;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        389: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        390: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        391: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        392: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        393: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        394: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        395: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        396: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        397: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        398: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        399: begin
          verilogPut_size_429 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_430 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_432 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_435 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_436 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_439 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_440 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_443 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_444 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_447 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        400: begin
          case (verilogPut_size_429)
            0: begin
              verilogPut_Key_449 <= verilogPut_Key_0_432;
              verilogPut_Data_451 <= verilogPut_Data_0_435;
            end
            1: begin
              verilogPut_Key_449 <= verilogPut_Key_1_436;
              verilogPut_Data_451 <= verilogPut_Data_1_439;
            end
            2: begin
              verilogPut_Key_449 <= verilogPut_Key_2_440;
              verilogPut_Data_451 <= verilogPut_Data_2_443;
            end
            3: begin
              verilogPut_Key_449 <= verilogPut_Key_3_444;
              verilogPut_Data_451 <= verilogPut_Data_3_447;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        401: begin
          verilogPut_childIndex_509 <= verilogPut_Data_451;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        402: begin
          verilogPut_index_455 <= verilogPut_childIndex_509;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        403: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_455;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_455;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_455;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_455;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_455;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_455;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_455;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_455;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_455;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_455;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        404: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        405: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        406: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        407: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        408: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        409: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        410: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        411: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        412: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        413: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        414: begin
          verilogPut_size_456 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_457 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_459 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_462 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_463 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_466 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_467 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_470 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_471 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_474 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        415: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        416: begin
          verilogPut_Key_0_486 <= verilogPut_Key_0_459;
          verilogPut_Data_0_489 <= verilogPut_Data_0_462;
          verilogPut_Key_1_490 <= verilogPut_Key_1_463;
          verilogPut_Data_1_493 <= verilogPut_Data_1_466;
          verilogPut_size_483 <= 2;
          verilogPut_Key_0_459 <= verilogPut_Key_2_467;
          verilogPut_Data_0_462 <= verilogPut_Data_2_470;
          verilogPut_Key_1_463 <= verilogPut_Key_3_471;
          verilogPut_Data_1_466 <= verilogPut_Data_3_474;
          verilogPut_size_456 <= 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        417: begin
          verilogPut_root_512 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        418: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_512;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        419: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        420: begin
          verilogPut_leftIndex_510 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        421: begin
          if (verilogPut_leftIndex_510 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_514 <= 1;
          verilogPut_isFree_515 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        422: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_leftIndex_510;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_leftIndex_510;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_514;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_leftIndex_510;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_515;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        423: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        424: begin
          verilogPut_next_513 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        425: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_512;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_513;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        426: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        427: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        428: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        429: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_leftIndex_510;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_483;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_leftIndex_510;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_486;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_leftIndex_510;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_489;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_leftIndex_510;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_490;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_leftIndex_510;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_493;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_leftIndex_510;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_494;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_leftIndex_510;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_497;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_leftIndex_510;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_498;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_leftIndex_510;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_501;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        430: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        431: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        432: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        433: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        434: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        435: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        436: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        437: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        438: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        439: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_childIndex_509;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_456;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_childIndex_509;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_459;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_childIndex_509;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_462;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_childIndex_509;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_463;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_childIndex_509;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_466;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_childIndex_509;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_467;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_childIndex_509;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_470;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_childIndex_509;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_471;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_childIndex_509;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_474;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        440: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        441: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        442: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        443: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        444: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        445: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        446: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        447: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        448: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        449: begin
          case (verilogPut_size_483)
            1: begin
              verilogPut_Key_503 <= verilogPut_Key_0_486;
              verilogPut_Data_505 <= verilogPut_Data_0_489;
            end
            2: begin
              verilogPut_Key_503 <= verilogPut_Key_1_490;
              verilogPut_Data_505 <= verilogPut_Data_1_493;
            end
            3: begin
              verilogPut_Key_503 <= verilogPut_Key_2_494;
              verilogPut_Data_505 <= verilogPut_Data_2_497;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        450: begin
          verilogPut_Key_476 <= verilogPut_Key_0_459;
          verilogPut_Data_478 <= verilogPut_Data_0_462;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        451: begin
          verilogPut_midKey_511 <= (verilogPut_Key_503 + verilogPut_Key_476) / 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        452: begin
          case (verilogPut_size_429)
            0: begin
              verilogPut_Key_0_432 <= verilogPut_midKey_511;
              verilogPut_Data_0_435 <= verilogPut_leftIndex_510;
            end
            1: begin
              verilogPut_Key_1_436 <= verilogPut_midKey_511;
              verilogPut_Data_1_439 <= verilogPut_leftIndex_510;
            end
            2: begin
              verilogPut_Key_2_440 <= verilogPut_midKey_511;
              verilogPut_Data_2_443 <= verilogPut_leftIndex_510;
            end
            3: begin
              verilogPut_Key_3_444 <= verilogPut_midKey_511;
              verilogPut_Data_3_447 <= verilogPut_leftIndex_510;
            end
          endcase
          verilogPut_size_429 <= verilogPut_size_429+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        453: begin
          case (verilogPut_size_429)
            0: begin
              verilogPut_Key_0_432 <= verilogPut_midKey_511;
              verilogPut_Data_0_435 <= verilogPut_childIndex_509;
            end
            1: begin
              verilogPut_Key_1_436 <= verilogPut_midKey_511;
              verilogPut_Data_1_439 <= verilogPut_childIndex_509;
            end
            2: begin
              verilogPut_Key_2_440 <= verilogPut_midKey_511;
              verilogPut_Data_2_443 <= verilogPut_childIndex_509;
            end
            3: begin
              verilogPut_Key_3_444 <= verilogPut_midKey_511;
              verilogPut_Data_3_447 <= verilogPut_childIndex_509;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        454: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_428;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_429;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_428;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_432;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_428;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_435;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_428;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_436;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_428;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_439;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_428;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_440;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_428;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_443;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_428;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_444;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_428;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_447;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        455: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        456: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        457: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        458: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        459: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        460: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        461: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        462: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        463: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        464: begin
          verilogPut_pc <= 465;
        end
        465: begin
          verilogPut_BtreeIndex_110 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        466: begin
          verilogPut_index_86 <= verilogPut_BtreeIndex_110;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        467: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_86;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_86;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_86;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_86;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_86;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_86;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_86;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_86;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_86;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_86;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        468: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        469: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        470: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        471: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        472: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        473: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        474: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        475: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        476: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        477: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        478: begin
          verilogPut_size_87 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_88 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_90 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_93 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_94 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_97 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_98 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_101 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_102 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_105 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        479: begin
          if (verilogPut_isLeaf_88 == 0) begin
            verilogPut_pc <= 486;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        480: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 == verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 == verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 == verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 == verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        481: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        482: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        483: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Key_107 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Key_107 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Key_107 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Key_107 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        484: begin
          verilogPut_pc <= 492;
        end
        485: begin
          verilogPut_pc <= 492;
        end
        486: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 <= verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 >  verilogPut_Key_0_90 && verilogPut_k_0 <= verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 >  verilogPut_Key_1_94 && verilogPut_k_0 <= verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 >  verilogPut_Key_2_98 && verilogPut_k_0 <= verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        487: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        488: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        489: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_FoundKey_108 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_FoundKey_108 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_FoundKey_108 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_FoundKey_108 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
            case (verilogPut_size_87)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        490: begin
          verilogPut_BtreeIndex_110 <= verilogPut_Data_109;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        491: begin
          verilogPut_pc <= 466;
        end
        492: begin
          if (verilogPut_Found_106 == 0) begin
            verilogPut_pc <= 495;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        493: begin
          if (verilogPut_StuckIndex_111 == verilogPut_size_87) begin
            verilogPut_size_87 <= verilogPut_size_87+1;
          end
          case (verilogPut_StuckIndex_111)
            0: begin
              verilogPut_Key_0_90 <= verilogPut_k_0;
              verilogPut_Data_0_93 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_94 <= verilogPut_k_0;
              verilogPut_Data_1_97 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_98 <= verilogPut_k_0;
              verilogPut_Data_2_101 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_102 <= verilogPut_k_0;
              verilogPut_Data_3_105 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        494: begin
          verilogPut_pc <= 506;
        end
        495: begin
          verilogPut_notFull_517 <= verilogPut_size_87< 4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        496: begin
          if (verilogPut_notFull_517 == 0) begin
            verilogPut_pc <= 505;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        497: begin
          verilogPut_KeyCompares_0_91 <= verilogPut_k_0 <= verilogPut_Key_0_90 && 0 < verilogPut_size_87;
          verilogPut_KeyCollapse_0_92 <= 0;
          verilogPut_KeyCompares_1_95 <= verilogPut_k_0 >  verilogPut_Key_0_90 && verilogPut_k_0 <= verilogPut_Key_1_94 && 1 < verilogPut_size_87;
          verilogPut_KeyCollapse_1_96 <= 1;
          verilogPut_KeyCompares_2_99 <= verilogPut_k_0 >  verilogPut_Key_1_94 && verilogPut_k_0 <= verilogPut_Key_2_98 && 2 < verilogPut_size_87;
          verilogPut_KeyCollapse_2_100 <= 2;
          verilogPut_KeyCompares_3_103 <= verilogPut_k_0 >  verilogPut_Key_2_98 && verilogPut_k_0 <= verilogPut_Key_3_102 && 3 < verilogPut_size_87;
          verilogPut_KeyCollapse_3_104 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        498: begin
          if (verilogPut_KeyCompares_1_95) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_1_96;
          end
          if (verilogPut_KeyCompares_3_103) begin
            verilogPut_KeyCompares_2_99 <= 1;
            verilogPut_KeyCollapse_2_100 <= verilogPut_KeyCollapse_3_104;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        499: begin
          if (verilogPut_KeyCompares_2_99) begin
            verilogPut_KeyCompares_0_91 <= 1;
            verilogPut_KeyCollapse_0_92 <= verilogPut_KeyCollapse_2_100;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        500: begin
          if (verilogPut_KeyCompares_0_91) begin
            verilogPut_Found_106 <= 1;
            case (verilogPut_KeyCollapse_0_92)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_FoundKey_108 <= verilogPut_Key_0_90;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_FoundKey_108 <= verilogPut_Key_1_94;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_FoundKey_108 <= verilogPut_Key_2_98;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_FoundKey_108 <= verilogPut_Key_3_102;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          else begin
            verilogPut_Found_106 <= 0;
            case (verilogPut_size_87)
              0: begin
                verilogPut_StuckIndex_111 <= 0;
                verilogPut_Data_109 <= verilogPut_Data_0_93;
              end
              1: begin
                verilogPut_StuckIndex_111 <= 1;
                verilogPut_Data_109 <= verilogPut_Data_1_97;
              end
              2: begin
                verilogPut_StuckIndex_111 <= 2;
                verilogPut_Data_109 <= verilogPut_Data_2_101;
              end
              3: begin
                verilogPut_StuckIndex_111 <= 3;
                verilogPut_Data_109 <= verilogPut_Data_3_105;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        501: begin
          verilogPut_size_87 <= verilogPut_size_87+1;
          if (3 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_3_102 <= verilogPut_Key_2_98;
            verilogPut_Data_3_105 <= verilogPut_Data_2_101;
          end
          if (2 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_2_98 <= verilogPut_Key_1_94;
            verilogPut_Data_2_101 <= verilogPut_Data_1_97;
          end
          if (1 > verilogPut_StuckIndex_111) begin
            verilogPut_Key_1_94 <= verilogPut_Key_0_90;
            verilogPut_Data_1_97 <= verilogPut_Data_0_93;
          end
          case (verilogPut_StuckIndex_111)
            0: begin
              verilogPut_Key_0_90 <= verilogPut_k_0;
              verilogPut_Data_0_93 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_94 <= verilogPut_k_0;
              verilogPut_Data_1_97 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_98 <= verilogPut_k_0;
              verilogPut_Data_2_101 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_102 <= verilogPut_k_0;
              verilogPut_Data_3_105 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        502: begin
          verilogPut_Found_106 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        503: begin
          verilogPut_pc <= verilogPut_pc + 1;
        end
        504: begin
          verilogPut_pc <= 506;
        end
        505: begin
          verilogPut_pc <= 516;
        end
        506: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_86;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_87;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_86;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_90;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_86;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_93;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_86;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_94;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_86;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_97;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_86;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_98;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_86;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_101;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_86;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_102;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_86;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_105;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        507: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        508: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        509: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        510: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        511: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        512: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        513: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        514: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        515: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        516: begin
          verilogPut_pc <= 671;
        end
        517: begin
          verilogPut_pc <= 671;
        end
        518: begin
          verilogPut_full_117 <= verilogPut_size_60>=3 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        519: begin
          if (verilogPut_full_117 == 0) begin
            verilogPut_pc <= 669;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        520: begin
          if (verilogPut_found_116 == 0) begin
            verilogPut_pc <= 594;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        521: begin
          verilogPut_index_518 <= verilogPut_parent_114;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        522: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_518;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_518;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_518;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_518;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_518;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_518;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_518;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_518;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_518;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_518;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        523: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        524: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        525: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        526: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        527: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        528: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        529: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        530: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        531: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        532: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        533: begin
          verilogPut_size_519 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_520 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_522 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_525 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_526 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_529 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_530 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_533 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_534 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_537 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        534: begin
          case (verilogPut_childInparent_115)
            0: begin
              verilogPut_childKey_626 <= verilogPut_Key_0_522;
              verilogPut_childData_627 <= verilogPut_Data_0_525;
            end
            1: begin
              verilogPut_childKey_626 <= verilogPut_Key_1_526;
              verilogPut_childData_627 <= verilogPut_Data_1_529;
            end
            2: begin
              verilogPut_childKey_626 <= verilogPut_Key_2_530;
              verilogPut_childData_627 <= verilogPut_Data_2_533;
            end
            3: begin
              verilogPut_childKey_626 <= verilogPut_Key_3_534;
              verilogPut_childData_627 <= verilogPut_Data_3_537;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        535: begin
          verilogPut_index_545 <= verilogPut_childData_627;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        536: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_545;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_545;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_545;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_545;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_545;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_545;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_545;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_545;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_545;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_545;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        537: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        538: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        539: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        540: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        541: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        542: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        543: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        544: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        545: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        546: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        547: begin
          verilogPut_size_546 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_547 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_549 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_552 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_553 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_556 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_557 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_560 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_561 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_564 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        548: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        549: begin
          verilogPut_Key_0_576 <= verilogPut_Key_0_549;
          verilogPut_Data_0_579 <= verilogPut_Data_0_552;
          verilogPut_size_573 <= 1;
          verilogPut_Data_1_583 <= verilogPut_Data_1_556;
          verilogPut_childKey_626 <= verilogPut_Key_1_553;
          verilogPut_Key_0_549 <= verilogPut_Key_2_557;
          verilogPut_Data_0_552 <= verilogPut_Data_2_560;
          verilogPut_Key_1_553 <= verilogPut_Key_3_561;
          verilogPut_Data_1_556 <= verilogPut_Data_3_564;
          verilogPut_size_546 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        550: begin
          verilogPut_root_631 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        551: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_631;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        552: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        553: begin
          verilogPut_indexLeft_628 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        554: begin
          if (verilogPut_indexLeft_628 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_633 <= 0;
          verilogPut_isFree_634 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        555: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexLeft_628;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexLeft_628;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_633;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_628;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_634;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        556: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        557: begin
          verilogPut_next_632 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        558: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_631;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_632;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        559: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        560: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        561: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        562: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexLeft_628;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_573;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexLeft_628;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_576;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexLeft_628;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_579;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexLeft_628;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_580;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexLeft_628;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_583;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexLeft_628;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_584;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexLeft_628;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_587;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexLeft_628;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_588;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexLeft_628;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_591;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        563: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        564: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        565: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        566: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        567: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        568: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        569: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        570: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        571: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        572: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_childData_627;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_546;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_childData_627;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_549;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_childData_627;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_552;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_childData_627;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_553;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_childData_627;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_556;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_childData_627;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_557;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_childData_627;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_560;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_childData_627;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_561;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_childData_627;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_564;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        573: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        574: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        575: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        576: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        577: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        578: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        579: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        580: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        581: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        582: begin
          verilogPut_size_519 <= verilogPut_size_519+1;
          if (3 > verilogPut_childInparent_115) begin
            verilogPut_Key_3_534 <= verilogPut_Key_2_530;
            verilogPut_Data_3_537 <= verilogPut_Data_2_533;
          end
          if (2 > verilogPut_childInparent_115) begin
            verilogPut_Key_2_530 <= verilogPut_Key_1_526;
            verilogPut_Data_2_533 <= verilogPut_Data_1_529;
          end
          if (1 > verilogPut_childInparent_115) begin
            verilogPut_Key_1_526 <= verilogPut_Key_0_522;
            verilogPut_Data_1_529 <= verilogPut_Data_0_525;
          end
          case (verilogPut_childInparent_115)
            0: begin
              verilogPut_Key_0_522 <= verilogPut_childKey_626;
              verilogPut_Data_0_525 <= verilogPut_indexLeft_628;
            end
            1: begin
              verilogPut_Key_1_526 <= verilogPut_childKey_626;
              verilogPut_Data_1_529 <= verilogPut_indexLeft_628;
            end
            2: begin
              verilogPut_Key_2_530 <= verilogPut_childKey_626;
              verilogPut_Data_2_533 <= verilogPut_indexLeft_628;
            end
            3: begin
              verilogPut_Key_3_534 <= verilogPut_childKey_626;
              verilogPut_Data_3_537 <= verilogPut_indexLeft_628;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        583: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_518;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_519;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_518;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_522;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_518;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_525;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_518;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_526;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_518;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_529;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_518;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_530;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_518;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_533;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_518;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_534;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_518;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_537;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        584: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        585: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        586: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        587: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        588: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        589: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        590: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        591: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        592: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        593: begin
          verilogPut_pc <= 668;
        end
        594: begin
          verilogPut_index_635 <= verilogPut_parent_114;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        595: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_635;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_635;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_635;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_635;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_635;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_635;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_635;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_635;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_635;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_635;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        596: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        597: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        598: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        599: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        600: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        601: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        602: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        603: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        604: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        605: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        606: begin
          verilogPut_size_636 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_637 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_639 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_642 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_643 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_646 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_647 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_650 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_651 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_654 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        607: begin
          case (verilogPut_size_636)
            0: begin
              verilogPut_Key_656 <= verilogPut_Key_0_639;
              verilogPut_Data_658 <= verilogPut_Data_0_642;
            end
            1: begin
              verilogPut_Key_656 <= verilogPut_Key_1_643;
              verilogPut_Data_658 <= verilogPut_Data_1_646;
            end
            2: begin
              verilogPut_Key_656 <= verilogPut_Key_2_647;
              verilogPut_Data_658 <= verilogPut_Data_2_650;
            end
            3: begin
              verilogPut_Key_656 <= verilogPut_Key_3_651;
              verilogPut_Data_658 <= verilogPut_Data_3_654;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        608: begin
          verilogPut_childData_744 <= verilogPut_Data_658;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        609: begin
          verilogPut_index_662 <= verilogPut_childData_744;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        610: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_662;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_662;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_662;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_662;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_662;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_662;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_662;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_662;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_662;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_662;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        611: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        612: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        613: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        614: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        615: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        616: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        617: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        618: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        619: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        620: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        621: begin
          verilogPut_size_663 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_664 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_666 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_669 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_670 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_673 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_674 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_677 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_678 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_681 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        622: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        623: begin
          verilogPut_Key_0_693 <= verilogPut_Key_0_666;
          verilogPut_Data_0_696 <= verilogPut_Data_0_669;
          verilogPut_size_690 <= 1;
          verilogPut_Data_1_700 <= verilogPut_Data_1_673;
          verilogPut_midKey_747 <= verilogPut_Key_1_670;
          verilogPut_Key_0_666 <= verilogPut_Key_2_674;
          verilogPut_Data_0_669 <= verilogPut_Data_2_677;
          verilogPut_Key_1_670 <= verilogPut_Key_3_678;
          verilogPut_Data_1_673 <= verilogPut_Data_3_681;
          verilogPut_size_663 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        624: begin
          verilogPut_root_748 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        625: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_748;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        626: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        627: begin
          verilogPut_indexLeft_745 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        628: begin
          if (verilogPut_indexLeft_745 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_750 <= 0;
          verilogPut_isFree_751 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        629: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_indexLeft_745;
          freeNext_21_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_indexLeft_745;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_750;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_745;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_751;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        630: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        631: begin
          verilogPut_next_749 <= freeNext_freeNext_21_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        632: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_root_748;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_749;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        633: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        634: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        635: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        636: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_indexLeft_745;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_690;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_indexLeft_745;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_693;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_indexLeft_745;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_696;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_indexLeft_745;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_697;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_indexLeft_745;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_700;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_indexLeft_745;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_701;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_indexLeft_745;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_704;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_indexLeft_745;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_705;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_indexLeft_745;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_708;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        637: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        638: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        639: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        640: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        641: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        642: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        643: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        644: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        645: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        646: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_childData_744;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_663;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_childData_744;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_666;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_childData_744;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_669;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_childData_744;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_670;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_childData_744;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_673;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_childData_744;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_674;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_childData_744;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_677;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_childData_744;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_678;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_childData_744;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_681;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        647: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        648: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        649: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        650: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        651: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        652: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        653: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        654: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        655: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        656: begin
          case (verilogPut_size_636)
            0: begin
              verilogPut_Key_0_639 <= verilogPut_midKey_747;
              verilogPut_Data_0_642 <= verilogPut_indexLeft_745;
            end
            1: begin
              verilogPut_Key_1_643 <= verilogPut_midKey_747;
              verilogPut_Data_1_646 <= verilogPut_indexLeft_745;
            end
            2: begin
              verilogPut_Key_2_647 <= verilogPut_midKey_747;
              verilogPut_Data_2_650 <= verilogPut_indexLeft_745;
            end
            3: begin
              verilogPut_Key_3_651 <= verilogPut_midKey_747;
              verilogPut_Data_3_654 <= verilogPut_indexLeft_745;
            end
          endcase
          verilogPut_size_636 <= verilogPut_size_636+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        657: begin
          case (verilogPut_size_636)
            0: begin
              verilogPut_Key_0_639 <= verilogPut_midKey_747;
              verilogPut_Data_0_642 <= verilogPut_childData_744;
            end
            1: begin
              verilogPut_Key_1_643 <= verilogPut_midKey_747;
              verilogPut_Data_1_646 <= verilogPut_childData_744;
            end
            2: begin
              verilogPut_Key_2_647 <= verilogPut_midKey_747;
              verilogPut_Data_2_650 <= verilogPut_childData_744;
            end
            3: begin
              verilogPut_Key_3_651 <= verilogPut_midKey_747;
              verilogPut_Data_3_654 <= verilogPut_childData_744;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        658: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_635;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_636;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_635;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_639;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_635;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_642;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_635;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_643;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_635;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_646;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_635;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_647;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_635;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_650;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_635;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_651;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_635;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_654;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        659: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        660: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        661: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        662: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        663: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        664: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        665: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        666: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        667: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        668: begin
          verilogPut_pc <= 670;
        end
        669: begin
          verilogPut_parent_114 <= verilogPut_child_113;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        670: begin
          verilogPut_pc <= 276;
        end
        671: begin
          verilogPut_position_779 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        672: begin
          verilogPut_index_752 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        673: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        674: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        675: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        676: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        677: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        678: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        679: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        680: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        681: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        682: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        683: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        684: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        685: begin
          if (verilogPut_isLeaf_754 == 0) begin
            verilogPut_pc <= 688;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        686: begin
          verilogPut_pc <= 1504;
        end
        687: begin
          verilogPut_pc <= 688;
        end
        688: begin
          verilogPut_success_869 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        689: begin
          verilogPut_index_783 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        690: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_783;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_783;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_783;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_783;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_783;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_783;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_783;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_783;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_783;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_783;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        691: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        692: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        693: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        694: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        695: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        696: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        697: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        698: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        699: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        700: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        701: begin
          verilogPut_size_784 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_785 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_787 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_790 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_791 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_794 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_795 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_798 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_799 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_802 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        702: begin
          verilogPut_test_870 <= verilogPut_size_784==1 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        703: begin
          if (verilogPut_test_870 == 0) begin
            verilogPut_pc <= 773;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        704: begin
          verilogPut_indexLeft_866 <= verilogPut_Data_0_790;
          verilogPut_indexRight_867 <= verilogPut_Data_1_794;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        705: begin
          verilogPut_index_810 <= verilogPut_indexLeft_866;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        706: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_810;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_810;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_810;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_810;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_810;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_810;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_810;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_810;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_810;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_810;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        707: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        708: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        709: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        710: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        711: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        712: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        713: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        714: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        715: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        716: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        717: begin
          verilogPut_size_811 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_812 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_814 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_817 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_818 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_821 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_822 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_825 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_826 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_829 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        718: begin
          verilogPut_index_837 <= verilogPut_indexRight_867;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        719: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_837;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_837;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_837;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_837;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_837;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_837;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_837;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_837;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_837;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_837;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        720: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        721: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        722: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        723: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        724: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        725: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        726: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        727: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        728: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        729: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        730: begin
          verilogPut_size_838 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_839 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_841 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_844 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_845 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_848 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_849 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_852 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_853 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_856 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        731: begin
          if (verilogPut_isLeaf_812 == 0) begin
            verilogPut_pc <= 773;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        732: begin
          if (verilogPut_isLeaf_839 == 0) begin
            verilogPut_pc <= 772;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        733: begin
          verilogPut_MergeSuccess_809 <= 0;
          case (verilogPut_size_811)
            0: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                4: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        734: begin
          if (verilogPut_MergeSuccess_809 == 0) begin
            verilogPut_pc <= 738;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        735: begin
          verilogPut_MergeSuccess_809 <= 0;
          case (verilogPut_size_784)
            0: begin
              case (verilogPut_size_811)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_814;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_817;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_814;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_817;
                  verilogPut_Key_1_791 <= verilogPut_Key_1_818;
                  verilogPut_Data_1_794 <= verilogPut_Data_1_821;
                  verilogPut_size_784 <= verilogPut_size_784 + 2;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_814;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_817;
                  verilogPut_Key_1_791 <= verilogPut_Key_1_818;
                  verilogPut_Data_1_794 <= verilogPut_Data_1_821;
                  verilogPut_Key_2_795 <= verilogPut_Key_2_822;
                  verilogPut_Data_2_798 <= verilogPut_Data_2_825;
                  verilogPut_size_784 <= verilogPut_size_784 + 3;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                4: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_814;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_817;
                  verilogPut_Key_1_791 <= verilogPut_Key_1_818;
                  verilogPut_Data_1_794 <= verilogPut_Data_1_821;
                  verilogPut_Key_2_795 <= verilogPut_Key_2_822;
                  verilogPut_Data_2_798 <= verilogPut_Data_2_825;
                  verilogPut_Key_3_799 <= verilogPut_Key_3_826;
                  verilogPut_Data_3_802 <= verilogPut_Data_3_829;
                  verilogPut_size_784 <= verilogPut_size_784 + 4;
                  verilogPut_MergeSuccess_809 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_811)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_1_791 <= verilogPut_Key_0_814;
                  verilogPut_Data_1_794 <= verilogPut_Data_0_817;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_Key_1_791 <= verilogPut_Key_0_814;
                  verilogPut_Data_1_794 <= verilogPut_Data_0_817;
                  verilogPut_Key_2_795 <= verilogPut_Key_1_818;
                  verilogPut_Data_2_798 <= verilogPut_Data_1_821;
                  verilogPut_size_784 <= verilogPut_size_784 + 2;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                  verilogPut_Key_1_791 <= verilogPut_Key_0_814;
                  verilogPut_Data_1_794 <= verilogPut_Data_0_817;
                  verilogPut_Key_2_795 <= verilogPut_Key_1_818;
                  verilogPut_Data_2_798 <= verilogPut_Data_1_821;
                  verilogPut_Key_3_799 <= verilogPut_Key_2_822;
                  verilogPut_Data_3_802 <= verilogPut_Data_2_825;
                  verilogPut_size_784 <= verilogPut_size_784 + 3;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_811)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_2_795 <= verilogPut_Key_0_814;
                  verilogPut_Data_2_798 <= verilogPut_Data_0_817;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_Key_2_795 <= verilogPut_Key_0_814;
                  verilogPut_Data_2_798 <= verilogPut_Data_0_817;
                  verilogPut_Key_3_799 <= verilogPut_Key_1_818;
                  verilogPut_Data_3_802 <= verilogPut_Data_1_821;
                  verilogPut_size_784 <= verilogPut_size_784 + 2;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_811)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_3_799 <= verilogPut_Key_0_814;
                  verilogPut_Data_3_802 <= verilogPut_Data_0_817;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_811)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        736: begin
          verilogPut_MergeSuccess_809 <= 0;
          case (verilogPut_size_784)
            0: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_841;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_844;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_841;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_844;
                  verilogPut_Key_1_791 <= verilogPut_Key_1_845;
                  verilogPut_Data_1_794 <= verilogPut_Data_1_848;
                  verilogPut_size_784 <= verilogPut_size_784 + 2;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_841;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_844;
                  verilogPut_Key_1_791 <= verilogPut_Key_1_845;
                  verilogPut_Data_1_794 <= verilogPut_Data_1_848;
                  verilogPut_Key_2_795 <= verilogPut_Key_2_849;
                  verilogPut_Data_2_798 <= verilogPut_Data_2_852;
                  verilogPut_size_784 <= verilogPut_size_784 + 3;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                4: begin
                  verilogPut_Key_0_787 <= verilogPut_Key_0_841;
                  verilogPut_Data_0_790 <= verilogPut_Data_0_844;
                  verilogPut_Key_1_791 <= verilogPut_Key_1_845;
                  verilogPut_Data_1_794 <= verilogPut_Data_1_848;
                  verilogPut_Key_2_795 <= verilogPut_Key_2_849;
                  verilogPut_Data_2_798 <= verilogPut_Data_2_852;
                  verilogPut_Key_3_799 <= verilogPut_Key_3_853;
                  verilogPut_Data_3_802 <= verilogPut_Data_3_856;
                  verilogPut_size_784 <= verilogPut_size_784 + 4;
                  verilogPut_MergeSuccess_809 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_1_791 <= verilogPut_Key_0_841;
                  verilogPut_Data_1_794 <= verilogPut_Data_0_844;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_Key_1_791 <= verilogPut_Key_0_841;
                  verilogPut_Data_1_794 <= verilogPut_Data_0_844;
                  verilogPut_Key_2_795 <= verilogPut_Key_1_845;
                  verilogPut_Data_2_798 <= verilogPut_Data_1_848;
                  verilogPut_size_784 <= verilogPut_size_784 + 2;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                  verilogPut_Key_1_791 <= verilogPut_Key_0_841;
                  verilogPut_Data_1_794 <= verilogPut_Data_0_844;
                  verilogPut_Key_2_795 <= verilogPut_Key_1_845;
                  verilogPut_Data_2_798 <= verilogPut_Data_1_848;
                  verilogPut_Key_3_799 <= verilogPut_Key_2_849;
                  verilogPut_Data_3_802 <= verilogPut_Data_2_852;
                  verilogPut_size_784 <= verilogPut_size_784 + 3;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_2_795 <= verilogPut_Key_0_841;
                  verilogPut_Data_2_798 <= verilogPut_Data_0_844;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                  verilogPut_Key_2_795 <= verilogPut_Key_0_841;
                  verilogPut_Data_2_798 <= verilogPut_Data_0_844;
                  verilogPut_Key_3_799 <= verilogPut_Key_1_845;
                  verilogPut_Data_3_802 <= verilogPut_Data_1_848;
                  verilogPut_size_784 <= verilogPut_size_784 + 2;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                  verilogPut_Key_3_799 <= verilogPut_Key_0_841;
                  verilogPut_Data_3_802 <= verilogPut_Data_0_844;
                  verilogPut_size_784 <= verilogPut_size_784 + 1;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_838)
                0: begin
                  verilogPut_size_784 <= verilogPut_size_784 + 0;
                  verilogPut_MergeSuccess_809 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        737: begin
          verilogPut_pc <= 738;
        end
        738: begin
          if (verilogPut_MergeSuccess_809 == 0) begin
            verilogPut_pc <= 771;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        739: begin
          verilogPut_isLeaf_785 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        740: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_783;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_784;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckIsLeaf_20_index_50 <= verilogPut_index_783;
          verilogPut_stuckIsLeaf_20_value_51 <= verilogPut_isLeaf_785;
          stuckIsLeaf_20_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_783;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_787;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_783;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_790;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_783;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_791;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_783;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_794;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_783;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_795;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_783;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_798;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_783;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_799;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_783;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_802;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        741: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        742: begin
          if ((stuckIsLeaf_20_requestedAt < stuckIsLeaf_20_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        743: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        744: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        745: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        746: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        747: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        748: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        749: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        750: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        751: begin
          verilogPut_root_872 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        752: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_872;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        753: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        754: begin
          verilogPut_next_871 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_872;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexLeft_866;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_873 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        755: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_866;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_873;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        756: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        757: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexLeft_866;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_871;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        758: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        759: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        760: begin
          verilogPut_root_875 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        761: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_875;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        762: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        763: begin
          verilogPut_next_874 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_875;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_867;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_876 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        764: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_867;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_876;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        765: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        766: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_867;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_874;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        767: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        768: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        769: begin
          verilogPut_success_869 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        770: begin
          verilogPut_pc <= 771;
        end
        771: begin
          verilogPut_pc <= 772;
        end
        772: begin
          verilogPut_pc <= 773;
        end
        773: begin
          if (verilogPut_success_869 == 0) begin
            verilogPut_pc <= 776;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        774: begin
          verilogPut_pc <= 1504;
        end
        775: begin
          verilogPut_pc <= 776;
        end
        776: begin
          verilogPut_index_877 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        777: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_877;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_877;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_877;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_877;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_877;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_877;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_877;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_877;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_877;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_877;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        778: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        779: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        780: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        781: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        782: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        783: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        784: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        785: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        786: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        787: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        788: begin
          verilogPut_size_878 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_879 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_881 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_884 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_885 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_888 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_889 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_892 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_893 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_896 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        789: begin
          verilogPut_success_965 <= 0;
          if (verilogPut_size_878 != 1) begin
            verilogPut_pc <= 853;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        790: begin
          verilogPut_midKey_964 <= verilogPut_Key_0_881;
          verilogPut_indexLeft_962 <= verilogPut_Data_0_884;
          verilogPut_indexRight_963 <= verilogPut_Data_1_888;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        791: begin
          if (verilogPut_isLeaf_906 == 0) begin
            verilogPut_pc <= 793;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        792: begin
          verilogPut_pc <= 853;
        end
        793: begin
          if (verilogPut_isLeaf_933 == 0) begin
            verilogPut_pc <= 795;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        794: begin
          verilogPut_pc <= 853;
        end
        795: begin
          verilogPut_index_904 <= verilogPut_indexLeft_962;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        796: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_904;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_904;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_904;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_904;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_904;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_904;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_904;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_904;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_904;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_904;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        797: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        798: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        799: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        800: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        801: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        802: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        803: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        804: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        805: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        806: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        807: begin
          verilogPut_size_905 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_906 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_908 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_911 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_912 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_915 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_916 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_919 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_920 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_923 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        808: begin
          verilogPut_index_931 <= verilogPut_indexRight_963;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        809: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_931;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_931;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_931;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_931;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_931;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_931;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_931;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_931;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_931;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_931;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        810: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        811: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        812: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        813: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        814: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        815: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        816: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        817: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        818: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        819: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        820: begin
          verilogPut_size_932 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_933 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_935 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_938 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_939 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_942 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_943 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_946 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_947 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_950 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        821: begin
          verilogPut_MergeSuccess_903 <= 0;
          case (verilogPut_size_905)
            0: begin
              case (verilogPut_size_932)
                0: begin
                  verilogPut_Key_0_881 <= verilogPut_midKey_964;
                  verilogPut_Data_0_884 <= verilogPut_Data_0_911;
                  verilogPut_Data_1_888 <= verilogPut_Data_0_938;
                  verilogPut_size_878 <= 1;
                  verilogPut_MergeSuccess_903 <= 1;
                end
                1: begin
                  verilogPut_Key_0_881 <= verilogPut_midKey_964;
                  verilogPut_Data_0_884 <= verilogPut_Data_0_911;
                  verilogPut_Key_1_885 <= verilogPut_Key_0_935;
                  verilogPut_Data_1_888 <= verilogPut_Data_0_938;
                  verilogPut_Data_2_892 <= verilogPut_Data_1_942;
                  verilogPut_size_878 <= 2;
                  verilogPut_MergeSuccess_903 <= 1;
                end
                2: begin
                  verilogPut_Key_0_881 <= verilogPut_midKey_964;
                  verilogPut_Data_0_884 <= verilogPut_Data_0_911;
                  verilogPut_Key_1_885 <= verilogPut_Key_0_935;
                  verilogPut_Data_1_888 <= verilogPut_Data_0_938;
                  verilogPut_Key_2_889 <= verilogPut_Key_1_939;
                  verilogPut_Data_2_892 <= verilogPut_Data_1_942;
                  verilogPut_Data_3_896 <= verilogPut_Data_2_946;
                  verilogPut_size_878 <= 3;
                  verilogPut_MergeSuccess_903 <= 1;
                end
                3: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_932)
                0: begin
                  verilogPut_Key_0_881 <= verilogPut_Key_0_908;
                  verilogPut_Data_0_884 <= verilogPut_Data_0_911;
                  verilogPut_Key_1_885 <= verilogPut_midKey_964;
                  verilogPut_Data_1_888 <= verilogPut_Data_1_915;
                  verilogPut_Data_2_892 <= verilogPut_Data_0_938;
                  verilogPut_size_878 <= 2;
                  verilogPut_MergeSuccess_903 <= 1;
                end
                1: begin
                  verilogPut_Key_0_881 <= verilogPut_Key_0_908;
                  verilogPut_Data_0_884 <= verilogPut_Data_0_911;
                  verilogPut_Key_1_885 <= verilogPut_midKey_964;
                  verilogPut_Data_1_888 <= verilogPut_Data_1_915;
                  verilogPut_Key_2_889 <= verilogPut_Key_0_935;
                  verilogPut_Data_2_892 <= verilogPut_Data_0_938;
                  verilogPut_Data_3_896 <= verilogPut_Data_1_942;
                  verilogPut_size_878 <= 3;
                  verilogPut_MergeSuccess_903 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_932)
                0: begin
                  verilogPut_Key_0_881 <= verilogPut_Key_0_908;
                  verilogPut_Data_0_884 <= verilogPut_Data_0_911;
                  verilogPut_Key_1_885 <= verilogPut_Key_1_912;
                  verilogPut_Data_1_888 <= verilogPut_Data_1_915;
                  verilogPut_Key_2_889 <= verilogPut_midKey_964;
                  verilogPut_Data_2_892 <= verilogPut_Data_2_919;
                  verilogPut_Data_3_896 <= verilogPut_Data_0_938;
                  verilogPut_size_878 <= 3;
                  verilogPut_MergeSuccess_903 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_932)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        822: begin
          if (verilogPut_MergeSuccess_903 == 0) begin
            verilogPut_pc <= 853;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        823: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_877;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_878;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_877;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_881;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_877;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_884;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_877;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_885;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_877;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_888;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_877;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_889;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_877;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_892;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_877;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_893;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_877;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_896;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        824: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        825: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        826: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        827: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        828: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        829: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        830: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        831: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        832: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        833: begin
          verilogPut_root_968 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        834: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_968;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        835: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        836: begin
          verilogPut_next_967 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_968;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexLeft_962;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_969 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        837: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexLeft_962;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_969;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        838: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        839: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexLeft_962;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_967;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        840: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        841: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        842: begin
          verilogPut_root_971 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        843: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_971;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        844: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        845: begin
          verilogPut_next_970 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_971;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_963;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_972 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        846: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_963;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_972;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        847: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        848: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_963;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_970;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        849: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        850: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        851: begin
          verilogPut_success_965 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        852: begin
          verilogPut_pc <= 853;
        end
        853: begin
          if (verilogPut_success_965 == 0) begin
            verilogPut_pc <= 868;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        854: begin
          verilogPut_index_752 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        855: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        856: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        857: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        858: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        859: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        860: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        861: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        862: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        863: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        864: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        865: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        866: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        867: begin
          verilogPut_pc <= 868;
        end
        868: begin
          verilogPut_success_1033 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        869: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 935;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        870: begin
          verilogPut_size_1028 <= verilogPut_size_753;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        871: begin
          case (verilogPut_size_1028)
            1: begin
              verilogPut_indexLeft_1030 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1031 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_indexLeft_1030 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1031 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_indexLeft_1030 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1031 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        872: begin
          verilogPut_index_973 <= verilogPut_indexLeft_1030;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        873: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_973;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_973;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_973;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_973;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_973;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_973;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_973;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_973;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_973;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_973;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        874: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        875: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        876: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        877: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        878: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        879: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        880: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        881: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        882: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        883: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        884: begin
          verilogPut_size_974 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_975 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_977 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_980 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_981 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_984 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_985 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_988 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_989 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_992 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        885: begin
          verilogPut_index_1000 <= verilogPut_indexRight_1031;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        886: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1000;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1000;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1000;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1000;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1000;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1000;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1000;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1000;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1000;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1000;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        887: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        888: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        889: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        890: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        891: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        892: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        893: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        894: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        895: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        896: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        897: begin
          verilogPut_size_1001 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1002 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1004 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1007 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1008 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1011 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1012 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1015 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1016 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1019 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        898: begin
          if (verilogPut_isLeaf_975 == 0) begin
            verilogPut_pc <= 935;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        899: begin
          if (verilogPut_isLeaf_1002 == 0) begin
            verilogPut_pc <= 934;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        900: begin
          verilogPut_MergeSuccess_999 <= 0;
          case (verilogPut_size_974)
            0: begin
              case (verilogPut_size_1001)
                0: begin
                  verilogPut_size_974 <= verilogPut_size_974 + 0;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                1: begin
                  verilogPut_Key_0_977 <= verilogPut_Key_0_1004;
                  verilogPut_Data_0_980 <= verilogPut_Data_0_1007;
                  verilogPut_size_974 <= verilogPut_size_974 + 1;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                2: begin
                  verilogPut_Key_0_977 <= verilogPut_Key_0_1004;
                  verilogPut_Data_0_980 <= verilogPut_Data_0_1007;
                  verilogPut_Key_1_981 <= verilogPut_Key_1_1008;
                  verilogPut_Data_1_984 <= verilogPut_Data_1_1011;
                  verilogPut_size_974 <= verilogPut_size_974 + 2;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                3: begin
                  verilogPut_Key_0_977 <= verilogPut_Key_0_1004;
                  verilogPut_Data_0_980 <= verilogPut_Data_0_1007;
                  verilogPut_Key_1_981 <= verilogPut_Key_1_1008;
                  verilogPut_Data_1_984 <= verilogPut_Data_1_1011;
                  verilogPut_Key_2_985 <= verilogPut_Key_2_1012;
                  verilogPut_Data_2_988 <= verilogPut_Data_2_1015;
                  verilogPut_size_974 <= verilogPut_size_974 + 3;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                4: begin
                  verilogPut_Key_0_977 <= verilogPut_Key_0_1004;
                  verilogPut_Data_0_980 <= verilogPut_Data_0_1007;
                  verilogPut_Key_1_981 <= verilogPut_Key_1_1008;
                  verilogPut_Data_1_984 <= verilogPut_Data_1_1011;
                  verilogPut_Key_2_985 <= verilogPut_Key_2_1012;
                  verilogPut_Data_2_988 <= verilogPut_Data_2_1015;
                  verilogPut_Key_3_989 <= verilogPut_Key_3_1016;
                  verilogPut_Data_3_992 <= verilogPut_Data_3_1019;
                  verilogPut_size_974 <= verilogPut_size_974 + 4;
                  verilogPut_MergeSuccess_999 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1001)
                0: begin
                  verilogPut_size_974 <= verilogPut_size_974 + 0;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                1: begin
                  verilogPut_Key_1_981 <= verilogPut_Key_0_1004;
                  verilogPut_Data_1_984 <= verilogPut_Data_0_1007;
                  verilogPut_size_974 <= verilogPut_size_974 + 1;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                2: begin
                  verilogPut_Key_1_981 <= verilogPut_Key_0_1004;
                  verilogPut_Data_1_984 <= verilogPut_Data_0_1007;
                  verilogPut_Key_2_985 <= verilogPut_Key_1_1008;
                  verilogPut_Data_2_988 <= verilogPut_Data_1_1011;
                  verilogPut_size_974 <= verilogPut_size_974 + 2;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                3: begin
                  verilogPut_Key_1_981 <= verilogPut_Key_0_1004;
                  verilogPut_Data_1_984 <= verilogPut_Data_0_1007;
                  verilogPut_Key_2_985 <= verilogPut_Key_1_1008;
                  verilogPut_Data_2_988 <= verilogPut_Data_1_1011;
                  verilogPut_Key_3_989 <= verilogPut_Key_2_1012;
                  verilogPut_Data_3_992 <= verilogPut_Data_2_1015;
                  verilogPut_size_974 <= verilogPut_size_974 + 3;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1001)
                0: begin
                  verilogPut_size_974 <= verilogPut_size_974 + 0;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                1: begin
                  verilogPut_Key_2_985 <= verilogPut_Key_0_1004;
                  verilogPut_Data_2_988 <= verilogPut_Data_0_1007;
                  verilogPut_size_974 <= verilogPut_size_974 + 1;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                2: begin
                  verilogPut_Key_2_985 <= verilogPut_Key_0_1004;
                  verilogPut_Data_2_988 <= verilogPut_Data_0_1007;
                  verilogPut_Key_3_989 <= verilogPut_Key_1_1008;
                  verilogPut_Data_3_992 <= verilogPut_Data_1_1011;
                  verilogPut_size_974 <= verilogPut_size_974 + 2;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1001)
                0: begin
                  verilogPut_size_974 <= verilogPut_size_974 + 0;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                1: begin
                  verilogPut_Key_3_989 <= verilogPut_Key_0_1004;
                  verilogPut_Data_3_992 <= verilogPut_Data_0_1007;
                  verilogPut_size_974 <= verilogPut_size_974 + 1;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1001)
                0: begin
                  verilogPut_size_974 <= verilogPut_size_974 + 0;
                  verilogPut_MergeSuccess_999 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        901: begin
          if (verilogPut_MergeSuccess_999 == 0) begin
            verilogPut_pc <= 933;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        902: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          verilogPut_success_1033 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        903: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_973;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_974;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_973;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_977;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_973;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_980;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_973;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_981;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_973;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_984;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_973;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_985;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_973;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_988;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_973;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_989;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_973;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_992;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        904: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        905: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        906: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        907: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        908: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        909: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        910: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        911: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        912: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        913: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        914: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        915: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        916: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        917: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        918: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        919: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        920: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        921: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        922: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        923: begin
          verilogPut_root_1036 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        924: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1036;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        925: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        926: begin
          verilogPut_next_1035 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1036;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1031;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1037 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        927: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1031;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1037;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        928: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        929: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1031;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1035;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        930: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        931: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        932: begin
          verilogPut_pc <= 933;
        end
        933: begin
          verilogPut_pc <= 934;
        end
        934: begin
          verilogPut_pc <= 935;
        end
        935: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1004;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        936: begin
          verilogPut_success_1098 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        937: begin
          verilogPut_size_1093 <= verilogPut_size_753;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        938: begin
          case (verilogPut_size_1093)
            1: begin
              verilogPut_indexLeft_1095 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1096 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_indexLeft_1095 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1096 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_indexLeft_1095 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1096 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        939: begin
          verilogPut_index_1038 <= verilogPut_indexLeft_1095;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        940: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1038;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1038;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1038;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1038;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1038;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1038;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1038;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1038;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1038;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1038;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        941: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        942: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        943: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        944: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        945: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        946: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        947: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        948: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        949: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        950: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        951: begin
          verilogPut_size_1039 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1040 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1042 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1045 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1046 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1049 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1050 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1053 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1054 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1057 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        952: begin
          verilogPut_index_1065 <= verilogPut_indexRight_1096;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        953: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1065;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1065;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1065;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1065;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1065;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1065;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1065;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1065;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1065;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1065;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        954: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        955: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        956: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        957: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        958: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        959: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        960: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        961: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        962: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        963: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        964: begin
          verilogPut_size_1066 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1067 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1069 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1072 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1073 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1076 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1077 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1080 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1081 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1084 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        965: begin
          if (verilogPut_isLeaf_1040 == 0) begin
            verilogPut_pc <= 967;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        966: begin
          verilogPut_pc <= 1004;
        end
        967: begin
          if (verilogPut_isLeaf_1067 == 0) begin
            verilogPut_pc <= 969;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        968: begin
          verilogPut_pc <= 1004;
        end
        969: begin
          case (verilogPut_size_753)
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            4: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_size_753 <= verilogPut_size_753-1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        970: begin
          verilogPut_MergeSuccess_1064 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        971: begin
          case (verilogPut_size_1039)
            0: begin
              case (verilogPut_size_1066)
                0: begin
                  verilogPut_Key_0_1042 <= verilogPut_Key_773;
                  verilogPut_Data_1_1049 <= verilogPut_Data_0_1072;
                  verilogPut_size_1039 <= verilogPut_size_1039 + 1;
                  verilogPut_MergeSuccess_1064 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1042 <= verilogPut_Key_773;
                  verilogPut_Key_1_1046 <= verilogPut_Key_0_1069;
                  verilogPut_Data_1_1049 <= verilogPut_Data_0_1072;
                  verilogPut_Data_2_1053 <= verilogPut_Data_1_1076;
                  verilogPut_size_1039 <= verilogPut_size_1039 + 2;
                  verilogPut_MergeSuccess_1064 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1042 <= verilogPut_Key_773;
                  verilogPut_Key_1_1046 <= verilogPut_Key_0_1069;
                  verilogPut_Data_1_1049 <= verilogPut_Data_0_1072;
                  verilogPut_Key_2_1050 <= verilogPut_Key_1_1073;
                  verilogPut_Data_2_1053 <= verilogPut_Data_1_1076;
                  verilogPut_Data_3_1057 <= verilogPut_Data_2_1080;
                  verilogPut_size_1039 <= verilogPut_size_1039 + 3;
                  verilogPut_MergeSuccess_1064 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1066)
                0: begin
                  verilogPut_Key_1_1046 <= verilogPut_Key_773;
                  verilogPut_Data_2_1053 <= verilogPut_Data_0_1072;
                  verilogPut_size_1039 <= verilogPut_size_1039 + 1;
                  verilogPut_MergeSuccess_1064 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1046 <= verilogPut_Key_773;
                  verilogPut_Key_2_1050 <= verilogPut_Key_0_1069;
                  verilogPut_Data_2_1053 <= verilogPut_Data_0_1072;
                  verilogPut_Data_3_1057 <= verilogPut_Data_1_1076;
                  verilogPut_size_1039 <= verilogPut_size_1039 + 2;
                  verilogPut_MergeSuccess_1064 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1066)
                0: begin
                  verilogPut_Key_2_1050 <= verilogPut_Key_773;
                  verilogPut_Data_3_1057 <= verilogPut_Data_0_1072;
                  verilogPut_size_1039 <= verilogPut_size_1039 + 1;
                  verilogPut_MergeSuccess_1064 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1066)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1066)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        972: begin
          if (verilogPut_MergeSuccess_1064 == 0) begin
            verilogPut_pc <= 1004;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        973: begin
          verilogPut_success_1098 <= 1;
          case (verilogPut_size_753)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1095;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1095;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1095;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1095;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        974: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1038;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1039;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1038;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1042;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1038;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1045;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1038;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1046;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1038;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1049;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1038;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1050;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1038;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1053;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1038;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1054;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1038;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1057;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        975: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        976: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        977: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        978: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        979: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        980: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        981: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        982: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        983: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        984: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        985: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        986: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        987: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        988: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        989: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        990: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        991: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        992: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        993: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        994: begin
          verilogPut_root_1101 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        995: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1101;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        996: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        997: begin
          verilogPut_next_1100 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1101;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1096;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1102 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        998: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1096;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1102;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        999: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1000: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1096;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1100;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1001: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1002: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1003: begin
          verilogPut_pc <= 1004;
        end
        1004: begin
          verilogPut_index_752 <= verilogPut_position_779;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1005: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1006: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1007: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1008: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1009: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1010: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1011: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1012: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1013: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1014: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1015: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1016: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1017: begin
          verilogPut_index_780 <= 2;
          verilogPut_within_781 <= verilogPut_size_753>=3 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1018: begin
          if (verilogPut_within_781 == 0) begin
            verilogPut_pc <= 1159;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1019: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1087;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        1020: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_indexLeft_1159 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1160 <= verilogPut_Data_1_763;
            end
            1: begin
              verilogPut_indexLeft_1159 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1160 <= verilogPut_Data_2_767;
            end
            2: begin
              verilogPut_indexLeft_1159 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1160 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1021: begin
          verilogPut_index_1103 <= verilogPut_indexLeft_1159;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1022: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1103;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1103;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1103;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1103;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1103;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1103;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1103;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1103;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1103;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1103;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1023: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1024: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1025: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1026: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1027: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1028: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1029: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1030: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1031: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1032: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1033: begin
          verilogPut_size_1104 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1105 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1107 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1110 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1111 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1114 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1115 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1118 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1119 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1122 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1034: begin
          verilogPut_index_1130 <= verilogPut_indexRight_1160;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1035: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1130;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1130;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1130;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1130;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1130;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1130;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1130;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1130;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1130;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1130;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1036: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1037: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1038: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1039: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1040: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1041: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1042: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1043: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1044: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1045: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1046: begin
          verilogPut_size_1131 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1132 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1134 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1137 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1138 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1141 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1142 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1145 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1146 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1149 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1047: begin
          if (verilogPut_isLeaf_1105 == 0) begin
            verilogPut_pc <= 1087;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1048: begin
          if (verilogPut_isLeaf_1132 == 0) begin
            verilogPut_pc <= 1086;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1049: begin
          verilogPut_MergeSuccess_1129 <= 0;
          case (verilogPut_size_1104)
            0: begin
              case (verilogPut_size_1131)
                0: begin
                  verilogPut_size_1104 <= verilogPut_size_1104 + 0;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1107 <= verilogPut_Key_0_1134;
                  verilogPut_Data_0_1110 <= verilogPut_Data_0_1137;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 1;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1107 <= verilogPut_Key_0_1134;
                  verilogPut_Data_0_1110 <= verilogPut_Data_0_1137;
                  verilogPut_Key_1_1111 <= verilogPut_Key_1_1138;
                  verilogPut_Data_1_1114 <= verilogPut_Data_1_1141;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 2;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                3: begin
                  verilogPut_Key_0_1107 <= verilogPut_Key_0_1134;
                  verilogPut_Data_0_1110 <= verilogPut_Data_0_1137;
                  verilogPut_Key_1_1111 <= verilogPut_Key_1_1138;
                  verilogPut_Data_1_1114 <= verilogPut_Data_1_1141;
                  verilogPut_Key_2_1115 <= verilogPut_Key_2_1142;
                  verilogPut_Data_2_1118 <= verilogPut_Data_2_1145;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 3;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                4: begin
                  verilogPut_Key_0_1107 <= verilogPut_Key_0_1134;
                  verilogPut_Data_0_1110 <= verilogPut_Data_0_1137;
                  verilogPut_Key_1_1111 <= verilogPut_Key_1_1138;
                  verilogPut_Data_1_1114 <= verilogPut_Data_1_1141;
                  verilogPut_Key_2_1115 <= verilogPut_Key_2_1142;
                  verilogPut_Data_2_1118 <= verilogPut_Data_2_1145;
                  verilogPut_Key_3_1119 <= verilogPut_Key_3_1146;
                  verilogPut_Data_3_1122 <= verilogPut_Data_3_1149;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 4;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1131)
                0: begin
                  verilogPut_size_1104 <= verilogPut_size_1104 + 0;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1111 <= verilogPut_Key_0_1134;
                  verilogPut_Data_1_1114 <= verilogPut_Data_0_1137;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 1;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                2: begin
                  verilogPut_Key_1_1111 <= verilogPut_Key_0_1134;
                  verilogPut_Data_1_1114 <= verilogPut_Data_0_1137;
                  verilogPut_Key_2_1115 <= verilogPut_Key_1_1138;
                  verilogPut_Data_2_1118 <= verilogPut_Data_1_1141;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 2;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                3: begin
                  verilogPut_Key_1_1111 <= verilogPut_Key_0_1134;
                  verilogPut_Data_1_1114 <= verilogPut_Data_0_1137;
                  verilogPut_Key_2_1115 <= verilogPut_Key_1_1138;
                  verilogPut_Data_2_1118 <= verilogPut_Data_1_1141;
                  verilogPut_Key_3_1119 <= verilogPut_Key_2_1142;
                  verilogPut_Data_3_1122 <= verilogPut_Data_2_1145;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 3;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1131)
                0: begin
                  verilogPut_size_1104 <= verilogPut_size_1104 + 0;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                1: begin
                  verilogPut_Key_2_1115 <= verilogPut_Key_0_1134;
                  verilogPut_Data_2_1118 <= verilogPut_Data_0_1137;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 1;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                2: begin
                  verilogPut_Key_2_1115 <= verilogPut_Key_0_1134;
                  verilogPut_Data_2_1118 <= verilogPut_Data_0_1137;
                  verilogPut_Key_3_1119 <= verilogPut_Key_1_1138;
                  verilogPut_Data_3_1122 <= verilogPut_Data_1_1141;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 2;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1131)
                0: begin
                  verilogPut_size_1104 <= verilogPut_size_1104 + 0;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                1: begin
                  verilogPut_Key_3_1119 <= verilogPut_Key_0_1134;
                  verilogPut_Data_3_1122 <= verilogPut_Data_0_1137;
                  verilogPut_size_1104 <= verilogPut_size_1104 + 1;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1131)
                0: begin
                  verilogPut_size_1104 <= verilogPut_size_1104 + 0;
                  verilogPut_MergeSuccess_1129 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1050: begin
          if (verilogPut_MergeSuccess_1129 == 0) begin
            verilogPut_pc <= 1085;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1051: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          if (0>= verilogPut_index_780) begin
            verilogPut_Key_0_756 <= verilogPut_Key_1_760;
            verilogPut_Data_0_759 <= verilogPut_Data_1_763;
          end
          if (1>= verilogPut_index_780) begin
            verilogPut_Key_1_760 <= verilogPut_Key_2_764;
            verilogPut_Data_1_763 <= verilogPut_Data_2_767;
          end
          if (2>= verilogPut_index_780) begin
            verilogPut_Key_2_764 <= verilogPut_Key_3_768;
            verilogPut_Data_2_767 <= verilogPut_Data_3_771;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1052: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1053: begin
          if (verilogPut_index_780 == verilogPut_size_753) begin
            verilogPut_size_753 <= verilogPut_size_753+1;
          end
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1159;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1159;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1159;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1159;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1054: begin
          verilogPut_success_1162 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1055: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1103;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1104;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1103;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1107;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1103;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1110;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1103;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1111;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1103;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1114;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1103;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1115;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1103;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1118;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1103;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1119;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1103;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1122;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1056: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1057: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1058: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1059: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1060: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1061: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1062: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1063: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1064: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1065: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1066: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1067: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1068: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1069: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1070: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1071: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1072: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1073: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1074: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1075: begin
          verilogPut_root_1165 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1076: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1165;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1077: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1078: begin
          verilogPut_next_1164 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1165;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1160;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1166 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1079: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1160;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1166;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1080: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1081: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1160;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1164;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1082: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1083: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1084: begin
          verilogPut_pc <= 1085;
        end
        1085: begin
          verilogPut_pc <= 1086;
        end
        1086: begin
          verilogPut_pc <= 1087;
        end
        1087: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1158;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        1088: begin
          verilogPut_success_1228 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1089: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_indexLeft_1225 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1226 <= verilogPut_Data_1_763;
            end
            1: begin
              verilogPut_indexLeft_1225 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1226 <= verilogPut_Data_2_767;
            end
            2: begin
              verilogPut_indexLeft_1225 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1226 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1090: begin
          verilogPut_index_1167 <= verilogPut_indexLeft_1225;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1091: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1167;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1167;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1167;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1167;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1167;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1167;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1167;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1167;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1167;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1167;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1092: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1093: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1094: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1095: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1096: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1097: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1098: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1099: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1100: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1101: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1102: begin
          verilogPut_size_1168 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1169 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1171 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1174 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1175 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1178 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1179 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1182 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1183 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1186 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1103: begin
          verilogPut_index_1194 <= verilogPut_indexRight_1226;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1104: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1194;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1194;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1194;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1194;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1194;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1194;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1194;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1194;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1194;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1194;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1105: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1106: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1107: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1108: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1109: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1110: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1111: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1112: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1113: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1114: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1115: begin
          verilogPut_size_1195 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1196 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1198 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1201 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1202 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1205 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1206 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1209 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1210 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1213 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1116: begin
          if (verilogPut_isLeaf_1169 == 0) begin
            verilogPut_pc <= 1118;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1117: begin
          verilogPut_pc <= 1158;
        end
        1118: begin
          if (verilogPut_isLeaf_1196 == 0) begin
            verilogPut_pc <= 1120;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1119: begin
          verilogPut_pc <= 1158;
        end
        1120: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_midKey_1227 <= verilogPut_Key_0_756;
            end
            1: begin
              verilogPut_midKey_1227 <= verilogPut_Key_1_760;
            end
            2: begin
              verilogPut_midKey_1227 <= verilogPut_Key_2_764;
            end
            3: begin
              verilogPut_midKey_1227 <= verilogPut_Key_3_768;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1121: begin
          verilogPut_MergeSuccess_1193 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1122: begin
          case (verilogPut_size_1168)
            0: begin
              case (verilogPut_size_1195)
                0: begin
                  verilogPut_Key_0_1171 <= verilogPut_midKey_1227;
                  verilogPut_Data_1_1178 <= verilogPut_Data_0_1201;
                  verilogPut_size_1168 <= verilogPut_size_1168 + 1;
                  verilogPut_MergeSuccess_1193 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1171 <= verilogPut_midKey_1227;
                  verilogPut_Key_1_1175 <= verilogPut_Key_0_1198;
                  verilogPut_Data_1_1178 <= verilogPut_Data_0_1201;
                  verilogPut_Data_2_1182 <= verilogPut_Data_1_1205;
                  verilogPut_size_1168 <= verilogPut_size_1168 + 2;
                  verilogPut_MergeSuccess_1193 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1171 <= verilogPut_midKey_1227;
                  verilogPut_Key_1_1175 <= verilogPut_Key_0_1198;
                  verilogPut_Data_1_1178 <= verilogPut_Data_0_1201;
                  verilogPut_Key_2_1179 <= verilogPut_Key_1_1202;
                  verilogPut_Data_2_1182 <= verilogPut_Data_1_1205;
                  verilogPut_Data_3_1186 <= verilogPut_Data_2_1209;
                  verilogPut_size_1168 <= verilogPut_size_1168 + 3;
                  verilogPut_MergeSuccess_1193 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1195)
                0: begin
                  verilogPut_Key_1_1175 <= verilogPut_midKey_1227;
                  verilogPut_Data_2_1182 <= verilogPut_Data_0_1201;
                  verilogPut_size_1168 <= verilogPut_size_1168 + 1;
                  verilogPut_MergeSuccess_1193 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1175 <= verilogPut_midKey_1227;
                  verilogPut_Key_2_1179 <= verilogPut_Key_0_1198;
                  verilogPut_Data_2_1182 <= verilogPut_Data_0_1201;
                  verilogPut_Data_3_1186 <= verilogPut_Data_1_1205;
                  verilogPut_size_1168 <= verilogPut_size_1168 + 2;
                  verilogPut_MergeSuccess_1193 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1195)
                0: begin
                  verilogPut_Key_2_1179 <= verilogPut_midKey_1227;
                  verilogPut_Data_3_1186 <= verilogPut_Data_0_1201;
                  verilogPut_size_1168 <= verilogPut_size_1168 + 1;
                  verilogPut_MergeSuccess_1193 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1195)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1195)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1123: begin
          if (verilogPut_MergeSuccess_1193 == 0) begin
            verilogPut_pc <= 1158;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1124: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          if (0>= verilogPut_index_780) begin
            verilogPut_Key_0_756 <= verilogPut_Key_1_760;
            verilogPut_Data_0_759 <= verilogPut_Data_1_763;
          end
          if (1>= verilogPut_index_780) begin
            verilogPut_Key_1_760 <= verilogPut_Key_2_764;
            verilogPut_Data_1_763 <= verilogPut_Data_2_767;
          end
          if (2>= verilogPut_index_780) begin
            verilogPut_Key_2_764 <= verilogPut_Key_3_768;
            verilogPut_Data_2_767 <= verilogPut_Data_3_771;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1125: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1126: begin
          if (verilogPut_index_780 == verilogPut_size_753) begin
            verilogPut_size_753 <= verilogPut_size_753+1;
          end
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1225;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1225;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1225;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1225;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1127: begin
          verilogPut_success_1228 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1128: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1167;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1168;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1167;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1171;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1167;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1174;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1167;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1175;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1167;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1178;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1167;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1179;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1167;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1182;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1167;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1183;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1167;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1186;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1129: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1130: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1131: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1132: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1133: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1134: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1135: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1136: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1137: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1138: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1139: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1140: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1141: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1142: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1143: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1144: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1145: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1146: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1147: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1148: begin
          verilogPut_root_1231 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1149: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1231;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1150: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1151: begin
          verilogPut_next_1230 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1231;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1226;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1232 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1152: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1226;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1232;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1153: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1154: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1226;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1230;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1155: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1156: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1157: begin
          verilogPut_pc <= 1158;
        end
        1158: begin
          verilogPut_pc <= 1159;
        end
        1159: begin
          verilogPut_index_752 <= verilogPut_position_779;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1160: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1161: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1162: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1163: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1164: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1165: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1166: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1167: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1168: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1169: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1170: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1171: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1172: begin
          verilogPut_index_780 <= 1;
          verilogPut_within_781 <= verilogPut_size_753>=2 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1173: begin
          if (verilogPut_within_781 == 0) begin
            verilogPut_pc <= 1314;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1174: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1242;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        1175: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_indexLeft_1289 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1290 <= verilogPut_Data_1_763;
            end
            1: begin
              verilogPut_indexLeft_1289 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1290 <= verilogPut_Data_2_767;
            end
            2: begin
              verilogPut_indexLeft_1289 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1290 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1176: begin
          verilogPut_index_1233 <= verilogPut_indexLeft_1289;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1177: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1233;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1233;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1233;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1233;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1233;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1233;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1233;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1233;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1233;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1233;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1178: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1179: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1180: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1181: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1182: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1183: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1184: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1185: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1186: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1187: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1188: begin
          verilogPut_size_1234 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1235 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1237 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1240 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1241 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1244 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1245 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1248 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1249 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1252 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1189: begin
          verilogPut_index_1260 <= verilogPut_indexRight_1290;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1190: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1260;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1260;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1260;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1260;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1260;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1260;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1260;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1260;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1260;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1260;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1191: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1192: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1193: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1194: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1195: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1196: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1197: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1198: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1199: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1200: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1201: begin
          verilogPut_size_1261 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1262 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1264 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1267 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1268 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1271 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1272 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1275 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1276 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1279 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1202: begin
          if (verilogPut_isLeaf_1235 == 0) begin
            verilogPut_pc <= 1242;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1203: begin
          if (verilogPut_isLeaf_1262 == 0) begin
            verilogPut_pc <= 1241;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1204: begin
          verilogPut_MergeSuccess_1259 <= 0;
          case (verilogPut_size_1234)
            0: begin
              case (verilogPut_size_1261)
                0: begin
                  verilogPut_size_1234 <= verilogPut_size_1234 + 0;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1237 <= verilogPut_Key_0_1264;
                  verilogPut_Data_0_1240 <= verilogPut_Data_0_1267;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 1;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1237 <= verilogPut_Key_0_1264;
                  verilogPut_Data_0_1240 <= verilogPut_Data_0_1267;
                  verilogPut_Key_1_1241 <= verilogPut_Key_1_1268;
                  verilogPut_Data_1_1244 <= verilogPut_Data_1_1271;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 2;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                3: begin
                  verilogPut_Key_0_1237 <= verilogPut_Key_0_1264;
                  verilogPut_Data_0_1240 <= verilogPut_Data_0_1267;
                  verilogPut_Key_1_1241 <= verilogPut_Key_1_1268;
                  verilogPut_Data_1_1244 <= verilogPut_Data_1_1271;
                  verilogPut_Key_2_1245 <= verilogPut_Key_2_1272;
                  verilogPut_Data_2_1248 <= verilogPut_Data_2_1275;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 3;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                4: begin
                  verilogPut_Key_0_1237 <= verilogPut_Key_0_1264;
                  verilogPut_Data_0_1240 <= verilogPut_Data_0_1267;
                  verilogPut_Key_1_1241 <= verilogPut_Key_1_1268;
                  verilogPut_Data_1_1244 <= verilogPut_Data_1_1271;
                  verilogPut_Key_2_1245 <= verilogPut_Key_2_1272;
                  verilogPut_Data_2_1248 <= verilogPut_Data_2_1275;
                  verilogPut_Key_3_1249 <= verilogPut_Key_3_1276;
                  verilogPut_Data_3_1252 <= verilogPut_Data_3_1279;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 4;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1261)
                0: begin
                  verilogPut_size_1234 <= verilogPut_size_1234 + 0;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1241 <= verilogPut_Key_0_1264;
                  verilogPut_Data_1_1244 <= verilogPut_Data_0_1267;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 1;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                2: begin
                  verilogPut_Key_1_1241 <= verilogPut_Key_0_1264;
                  verilogPut_Data_1_1244 <= verilogPut_Data_0_1267;
                  verilogPut_Key_2_1245 <= verilogPut_Key_1_1268;
                  verilogPut_Data_2_1248 <= verilogPut_Data_1_1271;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 2;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                3: begin
                  verilogPut_Key_1_1241 <= verilogPut_Key_0_1264;
                  verilogPut_Data_1_1244 <= verilogPut_Data_0_1267;
                  verilogPut_Key_2_1245 <= verilogPut_Key_1_1268;
                  verilogPut_Data_2_1248 <= verilogPut_Data_1_1271;
                  verilogPut_Key_3_1249 <= verilogPut_Key_2_1272;
                  verilogPut_Data_3_1252 <= verilogPut_Data_2_1275;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 3;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1261)
                0: begin
                  verilogPut_size_1234 <= verilogPut_size_1234 + 0;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                1: begin
                  verilogPut_Key_2_1245 <= verilogPut_Key_0_1264;
                  verilogPut_Data_2_1248 <= verilogPut_Data_0_1267;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 1;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                2: begin
                  verilogPut_Key_2_1245 <= verilogPut_Key_0_1264;
                  verilogPut_Data_2_1248 <= verilogPut_Data_0_1267;
                  verilogPut_Key_3_1249 <= verilogPut_Key_1_1268;
                  verilogPut_Data_3_1252 <= verilogPut_Data_1_1271;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 2;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1261)
                0: begin
                  verilogPut_size_1234 <= verilogPut_size_1234 + 0;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                1: begin
                  verilogPut_Key_3_1249 <= verilogPut_Key_0_1264;
                  verilogPut_Data_3_1252 <= verilogPut_Data_0_1267;
                  verilogPut_size_1234 <= verilogPut_size_1234 + 1;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1261)
                0: begin
                  verilogPut_size_1234 <= verilogPut_size_1234 + 0;
                  verilogPut_MergeSuccess_1259 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1205: begin
          if (verilogPut_MergeSuccess_1259 == 0) begin
            verilogPut_pc <= 1240;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1206: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          if (0>= verilogPut_index_780) begin
            verilogPut_Key_0_756 <= verilogPut_Key_1_760;
            verilogPut_Data_0_759 <= verilogPut_Data_1_763;
          end
          if (1>= verilogPut_index_780) begin
            verilogPut_Key_1_760 <= verilogPut_Key_2_764;
            verilogPut_Data_1_763 <= verilogPut_Data_2_767;
          end
          if (2>= verilogPut_index_780) begin
            verilogPut_Key_2_764 <= verilogPut_Key_3_768;
            verilogPut_Data_2_767 <= verilogPut_Data_3_771;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1207: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1208: begin
          if (verilogPut_index_780 == verilogPut_size_753) begin
            verilogPut_size_753 <= verilogPut_size_753+1;
          end
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1289;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1289;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1289;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1289;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1209: begin
          verilogPut_success_1292 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1210: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1233;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1234;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1233;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1237;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1233;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1240;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1233;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1241;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1233;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1244;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1233;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1245;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1233;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1248;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1233;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1249;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1233;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1252;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1211: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1212: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1213: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1214: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1215: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1216: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1217: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1218: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1219: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1220: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1221: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1222: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1223: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1224: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1225: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1226: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1227: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1228: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1229: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1230: begin
          verilogPut_root_1295 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1231: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1295;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1232: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1233: begin
          verilogPut_next_1294 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1295;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1290;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1296 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1234: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1290;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1296;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1235: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1236: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1290;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1294;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1237: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1238: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1239: begin
          verilogPut_pc <= 1240;
        end
        1240: begin
          verilogPut_pc <= 1241;
        end
        1241: begin
          verilogPut_pc <= 1242;
        end
        1242: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1313;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        1243: begin
          verilogPut_success_1358 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1244: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_indexLeft_1355 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1356 <= verilogPut_Data_1_763;
            end
            1: begin
              verilogPut_indexLeft_1355 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1356 <= verilogPut_Data_2_767;
            end
            2: begin
              verilogPut_indexLeft_1355 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1356 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1245: begin
          verilogPut_index_1297 <= verilogPut_indexLeft_1355;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1246: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1297;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1297;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1297;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1297;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1297;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1297;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1297;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1297;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1297;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1297;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1247: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1248: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1249: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1250: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1251: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1252: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1253: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1254: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1255: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1256: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1257: begin
          verilogPut_size_1298 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1299 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1301 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1304 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1305 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1308 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1309 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1312 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1313 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1316 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1258: begin
          verilogPut_index_1324 <= verilogPut_indexRight_1356;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1259: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1324;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1324;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1324;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1324;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1324;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1324;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1324;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1324;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1324;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1324;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1260: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1261: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1262: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1263: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1264: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1265: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1266: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1267: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1268: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1269: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1270: begin
          verilogPut_size_1325 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1326 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1328 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1331 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1332 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1335 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1336 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1339 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1340 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1343 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1271: begin
          if (verilogPut_isLeaf_1299 == 0) begin
            verilogPut_pc <= 1273;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1272: begin
          verilogPut_pc <= 1313;
        end
        1273: begin
          if (verilogPut_isLeaf_1326 == 0) begin
            verilogPut_pc <= 1275;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1274: begin
          verilogPut_pc <= 1313;
        end
        1275: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_midKey_1357 <= verilogPut_Key_0_756;
            end
            1: begin
              verilogPut_midKey_1357 <= verilogPut_Key_1_760;
            end
            2: begin
              verilogPut_midKey_1357 <= verilogPut_Key_2_764;
            end
            3: begin
              verilogPut_midKey_1357 <= verilogPut_Key_3_768;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1276: begin
          verilogPut_MergeSuccess_1323 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1277: begin
          case (verilogPut_size_1298)
            0: begin
              case (verilogPut_size_1325)
                0: begin
                  verilogPut_Key_0_1301 <= verilogPut_midKey_1357;
                  verilogPut_Data_1_1308 <= verilogPut_Data_0_1331;
                  verilogPut_size_1298 <= verilogPut_size_1298 + 1;
                  verilogPut_MergeSuccess_1323 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1301 <= verilogPut_midKey_1357;
                  verilogPut_Key_1_1305 <= verilogPut_Key_0_1328;
                  verilogPut_Data_1_1308 <= verilogPut_Data_0_1331;
                  verilogPut_Data_2_1312 <= verilogPut_Data_1_1335;
                  verilogPut_size_1298 <= verilogPut_size_1298 + 2;
                  verilogPut_MergeSuccess_1323 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1301 <= verilogPut_midKey_1357;
                  verilogPut_Key_1_1305 <= verilogPut_Key_0_1328;
                  verilogPut_Data_1_1308 <= verilogPut_Data_0_1331;
                  verilogPut_Key_2_1309 <= verilogPut_Key_1_1332;
                  verilogPut_Data_2_1312 <= verilogPut_Data_1_1335;
                  verilogPut_Data_3_1316 <= verilogPut_Data_2_1339;
                  verilogPut_size_1298 <= verilogPut_size_1298 + 3;
                  verilogPut_MergeSuccess_1323 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1325)
                0: begin
                  verilogPut_Key_1_1305 <= verilogPut_midKey_1357;
                  verilogPut_Data_2_1312 <= verilogPut_Data_0_1331;
                  verilogPut_size_1298 <= verilogPut_size_1298 + 1;
                  verilogPut_MergeSuccess_1323 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1305 <= verilogPut_midKey_1357;
                  verilogPut_Key_2_1309 <= verilogPut_Key_0_1328;
                  verilogPut_Data_2_1312 <= verilogPut_Data_0_1331;
                  verilogPut_Data_3_1316 <= verilogPut_Data_1_1335;
                  verilogPut_size_1298 <= verilogPut_size_1298 + 2;
                  verilogPut_MergeSuccess_1323 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1325)
                0: begin
                  verilogPut_Key_2_1309 <= verilogPut_midKey_1357;
                  verilogPut_Data_3_1316 <= verilogPut_Data_0_1331;
                  verilogPut_size_1298 <= verilogPut_size_1298 + 1;
                  verilogPut_MergeSuccess_1323 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1325)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1325)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1278: begin
          if (verilogPut_MergeSuccess_1323 == 0) begin
            verilogPut_pc <= 1313;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1279: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          if (0>= verilogPut_index_780) begin
            verilogPut_Key_0_756 <= verilogPut_Key_1_760;
            verilogPut_Data_0_759 <= verilogPut_Data_1_763;
          end
          if (1>= verilogPut_index_780) begin
            verilogPut_Key_1_760 <= verilogPut_Key_2_764;
            verilogPut_Data_1_763 <= verilogPut_Data_2_767;
          end
          if (2>= verilogPut_index_780) begin
            verilogPut_Key_2_764 <= verilogPut_Key_3_768;
            verilogPut_Data_2_767 <= verilogPut_Data_3_771;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1280: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1281: begin
          if (verilogPut_index_780 == verilogPut_size_753) begin
            verilogPut_size_753 <= verilogPut_size_753+1;
          end
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1355;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1355;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1355;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1355;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1282: begin
          verilogPut_success_1358 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1283: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1297;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1298;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1297;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1301;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1297;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1304;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1297;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1305;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1297;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1308;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1297;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1309;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1297;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1312;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1297;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1313;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1297;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1316;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1284: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1285: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1286: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1287: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1288: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1289: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1290: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1291: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1292: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1293: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1294: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1295: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1296: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1297: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1298: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1299: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1300: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1301: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1302: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1303: begin
          verilogPut_root_1361 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1304: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1361;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1305: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1306: begin
          verilogPut_next_1360 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1361;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1356;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1362 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1307: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1356;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1362;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1308: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1309: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1356;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1360;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1310: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1311: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1312: begin
          verilogPut_pc <= 1313;
        end
        1313: begin
          verilogPut_pc <= 1314;
        end
        1314: begin
          verilogPut_index_752 <= verilogPut_position_779;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1315: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1316: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1317: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1318: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1319: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1320: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1321: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1322: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1323: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1324: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1325: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1326: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1327: begin
          verilogPut_index_780 <= 0;
          verilogPut_within_781 <= verilogPut_size_753>=1 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1328: begin
          if (verilogPut_within_781 == 0) begin
            verilogPut_pc <= 1469;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1329: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1397;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        1330: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_indexLeft_1419 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1420 <= verilogPut_Data_1_763;
            end
            1: begin
              verilogPut_indexLeft_1419 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1420 <= verilogPut_Data_2_767;
            end
            2: begin
              verilogPut_indexLeft_1419 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1420 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1331: begin
          verilogPut_index_1363 <= verilogPut_indexLeft_1419;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1332: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1363;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1363;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1363;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1363;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1363;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1363;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1363;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1363;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1363;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1363;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1333: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1334: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1335: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1336: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1337: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1338: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1339: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1340: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1341: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1342: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1343: begin
          verilogPut_size_1364 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1365 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1367 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1370 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1371 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1374 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1375 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1378 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1379 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1382 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1344: begin
          verilogPut_index_1390 <= verilogPut_indexRight_1420;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1345: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1390;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1390;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1390;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1390;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1390;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1390;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1390;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1390;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1390;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1390;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1346: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1347: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1348: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1349: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1350: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1351: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1352: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1353: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1354: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1355: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1356: begin
          verilogPut_size_1391 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1392 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1394 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1397 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1398 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1401 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1402 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1405 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1406 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1409 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1357: begin
          if (verilogPut_isLeaf_1365 == 0) begin
            verilogPut_pc <= 1397;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1358: begin
          if (verilogPut_isLeaf_1392 == 0) begin
            verilogPut_pc <= 1396;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1359: begin
          verilogPut_MergeSuccess_1389 <= 0;
          case (verilogPut_size_1364)
            0: begin
              case (verilogPut_size_1391)
                0: begin
                  verilogPut_size_1364 <= verilogPut_size_1364 + 0;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1367 <= verilogPut_Key_0_1394;
                  verilogPut_Data_0_1370 <= verilogPut_Data_0_1397;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 1;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1367 <= verilogPut_Key_0_1394;
                  verilogPut_Data_0_1370 <= verilogPut_Data_0_1397;
                  verilogPut_Key_1_1371 <= verilogPut_Key_1_1398;
                  verilogPut_Data_1_1374 <= verilogPut_Data_1_1401;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 2;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                3: begin
                  verilogPut_Key_0_1367 <= verilogPut_Key_0_1394;
                  verilogPut_Data_0_1370 <= verilogPut_Data_0_1397;
                  verilogPut_Key_1_1371 <= verilogPut_Key_1_1398;
                  verilogPut_Data_1_1374 <= verilogPut_Data_1_1401;
                  verilogPut_Key_2_1375 <= verilogPut_Key_2_1402;
                  verilogPut_Data_2_1378 <= verilogPut_Data_2_1405;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 3;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                4: begin
                  verilogPut_Key_0_1367 <= verilogPut_Key_0_1394;
                  verilogPut_Data_0_1370 <= verilogPut_Data_0_1397;
                  verilogPut_Key_1_1371 <= verilogPut_Key_1_1398;
                  verilogPut_Data_1_1374 <= verilogPut_Data_1_1401;
                  verilogPut_Key_2_1375 <= verilogPut_Key_2_1402;
                  verilogPut_Data_2_1378 <= verilogPut_Data_2_1405;
                  verilogPut_Key_3_1379 <= verilogPut_Key_3_1406;
                  verilogPut_Data_3_1382 <= verilogPut_Data_3_1409;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 4;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1391)
                0: begin
                  verilogPut_size_1364 <= verilogPut_size_1364 + 0;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1371 <= verilogPut_Key_0_1394;
                  verilogPut_Data_1_1374 <= verilogPut_Data_0_1397;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 1;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                2: begin
                  verilogPut_Key_1_1371 <= verilogPut_Key_0_1394;
                  verilogPut_Data_1_1374 <= verilogPut_Data_0_1397;
                  verilogPut_Key_2_1375 <= verilogPut_Key_1_1398;
                  verilogPut_Data_2_1378 <= verilogPut_Data_1_1401;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 2;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                3: begin
                  verilogPut_Key_1_1371 <= verilogPut_Key_0_1394;
                  verilogPut_Data_1_1374 <= verilogPut_Data_0_1397;
                  verilogPut_Key_2_1375 <= verilogPut_Key_1_1398;
                  verilogPut_Data_2_1378 <= verilogPut_Data_1_1401;
                  verilogPut_Key_3_1379 <= verilogPut_Key_2_1402;
                  verilogPut_Data_3_1382 <= verilogPut_Data_2_1405;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 3;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1391)
                0: begin
                  verilogPut_size_1364 <= verilogPut_size_1364 + 0;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                1: begin
                  verilogPut_Key_2_1375 <= verilogPut_Key_0_1394;
                  verilogPut_Data_2_1378 <= verilogPut_Data_0_1397;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 1;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                2: begin
                  verilogPut_Key_2_1375 <= verilogPut_Key_0_1394;
                  verilogPut_Data_2_1378 <= verilogPut_Data_0_1397;
                  verilogPut_Key_3_1379 <= verilogPut_Key_1_1398;
                  verilogPut_Data_3_1382 <= verilogPut_Data_1_1401;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 2;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1391)
                0: begin
                  verilogPut_size_1364 <= verilogPut_size_1364 + 0;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                1: begin
                  verilogPut_Key_3_1379 <= verilogPut_Key_0_1394;
                  verilogPut_Data_3_1382 <= verilogPut_Data_0_1397;
                  verilogPut_size_1364 <= verilogPut_size_1364 + 1;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1391)
                0: begin
                  verilogPut_size_1364 <= verilogPut_size_1364 + 0;
                  verilogPut_MergeSuccess_1389 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1360: begin
          if (verilogPut_MergeSuccess_1389 == 0) begin
            verilogPut_pc <= 1395;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1361: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          if (0>= verilogPut_index_780) begin
            verilogPut_Key_0_756 <= verilogPut_Key_1_760;
            verilogPut_Data_0_759 <= verilogPut_Data_1_763;
          end
          if (1>= verilogPut_index_780) begin
            verilogPut_Key_1_760 <= verilogPut_Key_2_764;
            verilogPut_Data_1_763 <= verilogPut_Data_2_767;
          end
          if (2>= verilogPut_index_780) begin
            verilogPut_Key_2_764 <= verilogPut_Key_3_768;
            verilogPut_Data_2_767 <= verilogPut_Data_3_771;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1362: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1363: begin
          if (verilogPut_index_780 == verilogPut_size_753) begin
            verilogPut_size_753 <= verilogPut_size_753+1;
          end
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1419;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1419;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1419;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1419;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1364: begin
          verilogPut_success_1422 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1365: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1363;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1364;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1363;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1367;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1363;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1370;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1363;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1371;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1363;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1374;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1363;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1375;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1363;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1378;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1363;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1379;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1363;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1382;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1366: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1367: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1368: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1369: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1370: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1371: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1372: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1373: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1374: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1375: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1376: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1377: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1378: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1379: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1380: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1381: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1382: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1383: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1384: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1385: begin
          verilogPut_root_1425 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1386: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1425;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1387: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1388: begin
          verilogPut_next_1424 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1425;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1420;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1426 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1389: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1420;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1426;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1390: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1391: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1420;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1424;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1392: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1393: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1394: begin
          verilogPut_pc <= 1395;
        end
        1395: begin
          verilogPut_pc <= 1396;
        end
        1396: begin
          verilogPut_pc <= 1397;
        end
        1397: begin
          if (verilogPut_position_779 == 0 && verilogPut_size_753 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_779 == 0 || verilogPut_size_753 < 1) begin
              verilogPut_pc <= 1468;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        1398: begin
          verilogPut_success_1488 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1399: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_indexLeft_1485 <= verilogPut_Data_0_759;
              verilogPut_indexRight_1486 <= verilogPut_Data_1_763;
            end
            1: begin
              verilogPut_indexLeft_1485 <= verilogPut_Data_1_763;
              verilogPut_indexRight_1486 <= verilogPut_Data_2_767;
            end
            2: begin
              verilogPut_indexLeft_1485 <= verilogPut_Data_2_767;
              verilogPut_indexRight_1486 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1400: begin
          verilogPut_index_1427 <= verilogPut_indexLeft_1485;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1401: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1427;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1427;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1427;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1427;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1427;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1427;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1427;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1427;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1427;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1427;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1402: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1403: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1404: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1405: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1406: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1407: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1408: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1409: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1410: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1411: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1412: begin
          verilogPut_size_1428 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1429 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1431 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1434 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1435 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1438 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1439 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1442 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1443 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1446 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1413: begin
          verilogPut_index_1454 <= verilogPut_indexRight_1486;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1414: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_1454;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_1454;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_1454;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_1454;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_1454;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_1454;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_1454;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_1454;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_1454;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_1454;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1415: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1416: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1417: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1418: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1419: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1420: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1421: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1422: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1423: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1424: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1425: begin
          verilogPut_size_1455 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_1456 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_1458 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_1461 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_1462 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_1465 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_1466 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_1469 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_1470 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_1473 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1426: begin
          if (verilogPut_isLeaf_1429 == 0) begin
            verilogPut_pc <= 1428;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1427: begin
          verilogPut_pc <= 1468;
        end
        1428: begin
          if (verilogPut_isLeaf_1456 == 0) begin
            verilogPut_pc <= 1430;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1429: begin
          verilogPut_pc <= 1468;
        end
        1430: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_midKey_1487 <= verilogPut_Key_0_756;
            end
            1: begin
              verilogPut_midKey_1487 <= verilogPut_Key_1_760;
            end
            2: begin
              verilogPut_midKey_1487 <= verilogPut_Key_2_764;
            end
            3: begin
              verilogPut_midKey_1487 <= verilogPut_Key_3_768;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1431: begin
          verilogPut_MergeSuccess_1453 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1432: begin
          case (verilogPut_size_1428)
            0: begin
              case (verilogPut_size_1455)
                0: begin
                  verilogPut_Key_0_1431 <= verilogPut_midKey_1487;
                  verilogPut_Data_1_1438 <= verilogPut_Data_0_1461;
                  verilogPut_size_1428 <= verilogPut_size_1428 + 1;
                  verilogPut_MergeSuccess_1453 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1431 <= verilogPut_midKey_1487;
                  verilogPut_Key_1_1435 <= verilogPut_Key_0_1458;
                  verilogPut_Data_1_1438 <= verilogPut_Data_0_1461;
                  verilogPut_Data_2_1442 <= verilogPut_Data_1_1465;
                  verilogPut_size_1428 <= verilogPut_size_1428 + 2;
                  verilogPut_MergeSuccess_1453 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1431 <= verilogPut_midKey_1487;
                  verilogPut_Key_1_1435 <= verilogPut_Key_0_1458;
                  verilogPut_Data_1_1438 <= verilogPut_Data_0_1461;
                  verilogPut_Key_2_1439 <= verilogPut_Key_1_1462;
                  verilogPut_Data_2_1442 <= verilogPut_Data_1_1465;
                  verilogPut_Data_3_1446 <= verilogPut_Data_2_1469;
                  verilogPut_size_1428 <= verilogPut_size_1428 + 3;
                  verilogPut_MergeSuccess_1453 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1455)
                0: begin
                  verilogPut_Key_1_1435 <= verilogPut_midKey_1487;
                  verilogPut_Data_2_1442 <= verilogPut_Data_0_1461;
                  verilogPut_size_1428 <= verilogPut_size_1428 + 1;
                  verilogPut_MergeSuccess_1453 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1435 <= verilogPut_midKey_1487;
                  verilogPut_Key_2_1439 <= verilogPut_Key_0_1458;
                  verilogPut_Data_2_1442 <= verilogPut_Data_0_1461;
                  verilogPut_Data_3_1446 <= verilogPut_Data_1_1465;
                  verilogPut_size_1428 <= verilogPut_size_1428 + 2;
                  verilogPut_MergeSuccess_1453 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1455)
                0: begin
                  verilogPut_Key_2_1439 <= verilogPut_midKey_1487;
                  verilogPut_Data_3_1446 <= verilogPut_Data_0_1461;
                  verilogPut_size_1428 <= verilogPut_size_1428 + 1;
                  verilogPut_MergeSuccess_1453 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1455)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1455)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1433: begin
          if (verilogPut_MergeSuccess_1453 == 0) begin
            verilogPut_pc <= 1468;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1434: begin
          verilogPut_size_753 <= verilogPut_size_753-1;
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          if (0>= verilogPut_index_780) begin
            verilogPut_Key_0_756 <= verilogPut_Key_1_760;
            verilogPut_Data_0_759 <= verilogPut_Data_1_763;
          end
          if (1>= verilogPut_index_780) begin
            verilogPut_Key_1_760 <= verilogPut_Key_2_764;
            verilogPut_Data_1_763 <= verilogPut_Data_2_767;
          end
          if (2>= verilogPut_index_780) begin
            verilogPut_Key_2_764 <= verilogPut_Key_3_768;
            verilogPut_Data_2_767 <= verilogPut_Data_3_771;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1435: begin
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_773 <= verilogPut_Key_0_756;
              verilogPut_Data_775 <= verilogPut_Data_0_759;
            end
            1: begin
              verilogPut_Key_773 <= verilogPut_Key_1_760;
              verilogPut_Data_775 <= verilogPut_Data_1_763;
            end
            2: begin
              verilogPut_Key_773 <= verilogPut_Key_2_764;
              verilogPut_Data_775 <= verilogPut_Data_2_767;
            end
            3: begin
              verilogPut_Key_773 <= verilogPut_Key_3_768;
              verilogPut_Data_775 <= verilogPut_Data_3_771;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1436: begin
          if (verilogPut_index_780 == verilogPut_size_753) begin
            verilogPut_size_753 <= verilogPut_size_753+1;
          end
          case (verilogPut_index_780)
            0: begin
              verilogPut_Key_0_756 <= verilogPut_Key_773;
              verilogPut_Data_0_759 <= verilogPut_indexLeft_1485;
            end
            1: begin
              verilogPut_Key_1_760 <= verilogPut_Key_773;
              verilogPut_Data_1_763 <= verilogPut_indexLeft_1485;
            end
            2: begin
              verilogPut_Key_2_764 <= verilogPut_Key_773;
              verilogPut_Data_2_767 <= verilogPut_indexLeft_1485;
            end
            3: begin
              verilogPut_Key_3_768 <= verilogPut_Key_773;
              verilogPut_Data_3_771 <= verilogPut_indexLeft_1485;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1437: begin
          verilogPut_success_1488 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1438: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_1427;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_1428;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_1427;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_1431;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_1427;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_1434;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_1427;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_1435;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_1427;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_1438;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_1427;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_1439;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_1427;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_1442;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_1427;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_1443;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_1427;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_1446;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1439: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1440: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1441: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1442: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1443: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1444: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1445: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1446: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1447: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1448: begin
          verilogPut_stuckSize_18_index_47 <= verilogPut_index_752;
          verilogPut_stuckSize_18_value_48 <= verilogPut_size_753;
          stuckSize_18_requestedAt <= step;
          verilogPut_stuckKeys_0_2_index_11 <= verilogPut_index_752;
          verilogPut_stuckKeys_0_2_value_12 <= verilogPut_Key_0_756;
          stuckKeys_0_2_requestedAt <= step;
          verilogPut_stuckData_0_4_index_14 <= verilogPut_index_752;
          verilogPut_stuckData_0_4_value_15 <= verilogPut_Data_0_759;
          stuckData_0_4_requestedAt <= step;
          verilogPut_stuckKeys_1_6_index_21 <= verilogPut_index_752;
          verilogPut_stuckKeys_1_6_value_22 <= verilogPut_Key_1_760;
          stuckKeys_1_6_requestedAt <= step;
          verilogPut_stuckData_1_8_index_24 <= verilogPut_index_752;
          verilogPut_stuckData_1_8_value_25 <= verilogPut_Data_1_763;
          stuckData_1_8_requestedAt <= step;
          verilogPut_stuckKeys_2_10_index_31 <= verilogPut_index_752;
          verilogPut_stuckKeys_2_10_value_32 <= verilogPut_Key_2_764;
          stuckKeys_2_10_requestedAt <= step;
          verilogPut_stuckData_2_12_index_34 <= verilogPut_index_752;
          verilogPut_stuckData_2_12_value_35 <= verilogPut_Data_2_767;
          stuckData_2_12_requestedAt <= step;
          verilogPut_stuckKeys_3_14_index_41 <= verilogPut_index_752;
          verilogPut_stuckKeys_3_14_value_42 <= verilogPut_Key_3_768;
          stuckKeys_3_14_requestedAt <= step;
          verilogPut_stuckData_3_16_index_44 <= verilogPut_index_752;
          verilogPut_stuckData_3_16_value_45 <= verilogPut_Data_3_771;
          stuckData_3_16_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1449: begin
          if ((stuckSize_18_requestedAt < stuckSize_18_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1450: begin
          if ((stuckKeys_0_2_requestedAt < stuckKeys_0_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1451: begin
          if ((stuckData_0_4_requestedAt < stuckData_0_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1452: begin
          if ((stuckKeys_1_6_requestedAt < stuckKeys_1_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1453: begin
          if ((stuckData_1_8_requestedAt < stuckData_1_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1454: begin
          if ((stuckKeys_2_10_requestedAt < stuckKeys_2_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1455: begin
          if ((stuckData_2_12_requestedAt < stuckData_2_12_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1456: begin
          if ((stuckKeys_3_14_requestedAt < stuckKeys_3_14_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1457: begin
          if ((stuckData_3_16_requestedAt < stuckData_3_16_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1458: begin
          verilogPut_root_1491 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1459: begin
          verilogPut_freeNext_21_index_204 <= verilogPut_root_1491;
          freeNext_21_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1460: begin
          if ((freeNext_21_requestedAt < freeNext_21_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1461: begin
          verilogPut_next_1490 <= freeNext_freeNext_21_result_0;
          verilogPut_freeNext_22_index_205 <= verilogPut_root_1491;
          verilogPut_freeNext_22_value_206 <= verilogPut_indexRight_1486;
          freeNext_22_requestedAt <= step;
          verilogPut_isFree_1492 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1462: begin
          verilogPut_stuckIsFree_23_index_207 <= verilogPut_indexRight_1486;
          verilogPut_stuckIsFree_23_value_208 <= verilogPut_isFree_1492;
          stuckIsFree_23_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1463: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1464: begin
          verilogPut_freeNext_22_index_205 <= verilogPut_indexRight_1486;
          verilogPut_freeNext_22_value_206 <= verilogPut_next_1490;
          freeNext_22_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1465: begin
          if ((freeNext_22_requestedAt < freeNext_22_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1466: begin
          if ((stuckIsFree_23_requestedAt < stuckIsFree_23_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1467: begin
          verilogPut_pc <= 1468;
        end
        1468: begin
          verilogPut_pc <= 1469;
        end
        1469: begin
          verilogPut_index_752 <= verilogPut_position_779;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1470: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1471: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1472: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1473: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1474: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1475: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1476: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1477: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1478: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1479: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1480: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1481: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1482: begin
          verilogPut_KeyCompares_0_757 <= verilogPut_k_0 <= verilogPut_Key_0_756 && 0 < verilogPut_size_753;
          verilogPut_KeyCollapse_0_758 <= 0;
          verilogPut_KeyCompares_1_761 <= verilogPut_k_0 >  verilogPut_Key_0_756 && verilogPut_k_0 <= verilogPut_Key_1_760 && 1 < verilogPut_size_753;
          verilogPut_KeyCollapse_1_762 <= 1;
          verilogPut_KeyCompares_2_765 <= verilogPut_k_0 >  verilogPut_Key_1_760 && verilogPut_k_0 <= verilogPut_Key_2_764 && 2 < verilogPut_size_753;
          verilogPut_KeyCollapse_2_766 <= 2;
          verilogPut_KeyCompares_3_769 <= verilogPut_k_0 >  verilogPut_Key_2_764 && verilogPut_k_0 <= verilogPut_Key_3_768 && 3 < verilogPut_size_753;
          verilogPut_KeyCollapse_3_770 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1483: begin
          if (verilogPut_KeyCompares_1_761) begin
            verilogPut_KeyCompares_0_757 <= 1;
            verilogPut_KeyCollapse_0_758 <= verilogPut_KeyCollapse_1_762;
          end
          if (verilogPut_KeyCompares_3_769) begin
            verilogPut_KeyCompares_2_765 <= 1;
            verilogPut_KeyCollapse_2_766 <= verilogPut_KeyCollapse_3_770;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1484: begin
          if (verilogPut_KeyCompares_2_765) begin
            verilogPut_KeyCompares_0_757 <= 1;
            verilogPut_KeyCollapse_0_758 <= verilogPut_KeyCollapse_2_766;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1485: begin
          if (verilogPut_KeyCompares_0_757) begin
            verilogPut_Found_772 <= 1;
            case (verilogPut_KeyCollapse_0_758)
              0: begin
                verilogPut_StuckIndex_777 <= 0;
                verilogPut_FoundKey_774 <= verilogPut_Key_0_756;
                verilogPut_Data_775 <= verilogPut_Data_0_759;
              end
              1: begin
                verilogPut_StuckIndex_777 <= 1;
                verilogPut_FoundKey_774 <= verilogPut_Key_1_760;
                verilogPut_Data_775 <= verilogPut_Data_1_763;
              end
              2: begin
                verilogPut_StuckIndex_777 <= 2;
                verilogPut_FoundKey_774 <= verilogPut_Key_2_764;
                verilogPut_Data_775 <= verilogPut_Data_2_767;
              end
              3: begin
                verilogPut_StuckIndex_777 <= 3;
                verilogPut_FoundKey_774 <= verilogPut_Key_3_768;
                verilogPut_Data_775 <= verilogPut_Data_3_771;
              end
            endcase
          end
          else begin
            verilogPut_Found_772 <= 0;
            case (verilogPut_size_753)
              0: begin
                verilogPut_StuckIndex_777 <= 0;
                verilogPut_Data_775 <= verilogPut_Data_0_759;
              end
              1: begin
                verilogPut_StuckIndex_777 <= 1;
                verilogPut_Data_775 <= verilogPut_Data_1_763;
              end
              2: begin
                verilogPut_StuckIndex_777 <= 2;
                verilogPut_Data_775 <= verilogPut_Data_2_767;
              end
              3: begin
                verilogPut_StuckIndex_777 <= 3;
                verilogPut_Data_775 <= verilogPut_Data_3_771;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1486: begin
          verilogPut_position_779 <= verilogPut_Data_775;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1487: begin
          verilogPut_index_752 <= verilogPut_position_779;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1488: begin
          verilogPut_stuckSize_17_index_46 <= verilogPut_index_752;
          stuckSize_17_requestedAt <= step;
          verilogPut_stuckIsLeaf_19_index_49 <= verilogPut_index_752;
          stuckIsLeaf_19_requestedAt <= step;
          verilogPut_stuckKeys_0_1_index_10 <= verilogPut_index_752;
          stuckKeys_0_1_requestedAt <= step;
          verilogPut_stuckData_0_3_index_13 <= verilogPut_index_752;
          stuckData_0_3_requestedAt <= step;
          verilogPut_stuckKeys_1_5_index_20 <= verilogPut_index_752;
          stuckKeys_1_5_requestedAt <= step;
          verilogPut_stuckData_1_7_index_23 <= verilogPut_index_752;
          stuckData_1_7_requestedAt <= step;
          verilogPut_stuckKeys_2_9_index_30 <= verilogPut_index_752;
          stuckKeys_2_9_requestedAt <= step;
          verilogPut_stuckData_2_11_index_33 <= verilogPut_index_752;
          stuckData_2_11_requestedAt <= step;
          verilogPut_stuckKeys_3_13_index_40 <= verilogPut_index_752;
          stuckKeys_3_13_requestedAt <= step;
          verilogPut_stuckData_3_15_index_43 <= verilogPut_index_752;
          stuckData_3_15_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1489: begin
          if ((stuckSize_17_requestedAt < stuckSize_17_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1490: begin
          if ((stuckIsLeaf_19_requestedAt < stuckIsLeaf_19_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1491: begin
          if ((stuckKeys_0_1_requestedAt < stuckKeys_0_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1492: begin
          if ((stuckData_0_3_requestedAt < stuckData_0_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1493: begin
          if ((stuckKeys_1_5_requestedAt < stuckKeys_1_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1494: begin
          if ((stuckData_1_7_requestedAt < stuckData_1_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1495: begin
          if ((stuckKeys_2_9_requestedAt < stuckKeys_2_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1496: begin
          if ((stuckData_2_11_requestedAt < stuckData_2_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1497: begin
          if ((stuckKeys_3_13_requestedAt < stuckKeys_3_13_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1498: begin
          if ((stuckData_3_15_requestedAt < stuckData_3_15_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1499: begin
          verilogPut_size_753 <= stuckSize_stuckSize_17_result_0;
          verilogPut_isLeaf_754 <= stuckIsLeaf_stuckIsLeaf_19_result_0;
          verilogPut_Key_0_756 <= stuckKeys_0_stuckKeys_0_1_result_0;
          verilogPut_Data_0_759 <= stuckData_0_stuckData_0_3_result_0;
          verilogPut_Key_1_760 <= stuckKeys_1_stuckKeys_1_5_result_0;
          verilogPut_Data_1_763 <= stuckData_1_stuckData_1_7_result_0;
          verilogPut_Key_2_764 <= stuckKeys_2_stuckKeys_2_9_result_0;
          verilogPut_Data_2_767 <= stuckData_2_stuckData_2_11_result_0;
          verilogPut_Key_3_768 <= stuckKeys_3_stuckKeys_3_13_result_0;
          verilogPut_Data_3_771 <= stuckData_3_stuckData_3_15_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1500: begin
          if (verilogPut_isLeaf_754 == 0) begin
            verilogPut_pc <= 1503;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        1501: begin
          verilogPut_pc <= 1504;
        end
        1502: begin
          verilogPut_pc <= 1504;
        end
        1503: begin
          verilogPut_pc <= 868;
        end
        default: verilogPut_stop <= 1;
      endcase
    end
  end
endmodule
