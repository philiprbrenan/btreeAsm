//-----------------------------------------------------------------------------
// Database on a chip test bench
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree;                                                                      // Test bench for database on a chip
  reg                    stop;                                                  // Program has stopped when this goes high
  reg                   clock;                                                  // Clock
  integer                step;                                                  // Step of the simulation
  integer            maxSteps;                                                  // Maximum number of steps to execute
  integer          returnCode;                                                  // Return code
  integer      processCurrent;                                                  // To ensure we get the same results in Java and Verilog we have to run the processes single threaded in a constant order

  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_stop||stuckData_stop||findAndInsert_stop;                                                             // Or of process stop fields

  initial begin
    returnCode = 0;
    maxSteps = 2000;
    for(step = -1; step < 0 || step < maxSteps && !stop; step = step + 1) begin // Steps below zero are run unconditionally to initialize each process so that Java and Verilog start in sync at step zero

      processCurrent = 0; clock = 0; #1; clock = 1; #1; // process_stuckIsLeaf_0000
      processCurrent = 1; clock = 0; #1; clock = 1; #1; // process_stuckIsFree_0001
      processCurrent = 2; clock = 0; #1; clock = 1; #1; // process_freeNext_0002
      processCurrent = 3; clock = 0; #1; clock = 1; #1; // process_stuckSize_0003
      processCurrent = 4; clock = 0; #1; clock = 1; #1; // process_stuckKeys_0004
      processCurrent = 5; clock = 0; #1; clock = 1; #1; // process_stuckData_0005
      processCurrent = 6; clock = 0; #1; clock = 1; #1; // process_findAndInsert_0006
      if (step >= 0) chipPrint();                                            // Steps prior to zero are for initialization to make Java and Verilog match
    end
    if (!stop) $finish(1); else $finish(0);                                // Set return code depending on whether the simulation halted
  end
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[32*1];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_7_result_0;
  integer stuckIsLeaf_7_requestedAt;
  integer stuckIsLeaf_7_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_7_returnCode;
  integer stuckIsLeaf_8_requestedAt;
  integer stuckIsLeaf_8_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_8_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_7_result_0 <= 0;
      stuckIsLeaf_7_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_7_returnCode <= 0;
      stuckIsLeaf_8_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_8_returnCode <= 0;
      stuckIsLeaf_memory[0] <= 1;
      stuckIsLeaf_memory[1] <= 0;
      stuckIsLeaf_memory[2] <= 0;
      stuckIsLeaf_memory[3] <= 0;
      stuckIsLeaf_memory[4] <= 0;
      stuckIsLeaf_memory[5] <= 0;
      stuckIsLeaf_memory[6] <= 0;
      stuckIsLeaf_memory[7] <= 0;
      stuckIsLeaf_memory[8] <= 0;
      stuckIsLeaf_memory[9] <= 0;
      stuckIsLeaf_memory[10] <= 0;
      stuckIsLeaf_memory[11] <= 0;
      stuckIsLeaf_memory[12] <= 0;
      stuckIsLeaf_memory[13] <= 0;
      stuckIsLeaf_memory[14] <= 0;
      stuckIsLeaf_memory[15] <= 0;
      stuckIsLeaf_memory[16] <= 0;
      stuckIsLeaf_memory[17] <= 0;
      stuckIsLeaf_memory[18] <= 0;
      stuckIsLeaf_memory[19] <= 0;
      stuckIsLeaf_memory[20] <= 0;
      stuckIsLeaf_memory[21] <= 0;
      stuckIsLeaf_memory[22] <= 0;
      stuckIsLeaf_memory[23] <= 0;
      stuckIsLeaf_memory[24] <= 0;
      stuckIsLeaf_memory[25] <= 0;
      stuckIsLeaf_memory[26] <= 0;
      stuckIsLeaf_memory[27] <= 0;
      stuckIsLeaf_memory[28] <= 0;
      stuckIsLeaf_memory[29] <= 0;
      stuckIsLeaf_memory[30] <= 0;
      stuckIsLeaf_memory[31] <= 0;
    end
    else if (processCurrent == 0) begin
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_7_result_0 <= stuckIsLeaf_memory[findAndInsert_stuckIsLeaf_7_index_35*1+0];
            stuckIsLeaf_7_finishedAt <= step;
          end
          else if ((stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step)) begin
            stuckIsLeaf_memory[findAndInsert_stuckIsLeaf_8_index_36*1+0] <= findAndInsert_stuckIsLeaf_8_value_37;
            stuckIsLeaf_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[32*1];
  integer stuckIsFree_11_requestedAt;
  integer stuckIsFree_11_finishedAt;
  integer stuckIsFree_stuckIsFree_11_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_11_finishedAt <= -1;
      stuckIsFree_stuckIsFree_11_returnCode <= 0;
      stuckIsFree_memory[0] <= 0;
      stuckIsFree_memory[1] <= 1;
      stuckIsFree_memory[2] <= 1;
      stuckIsFree_memory[3] <= 1;
      stuckIsFree_memory[4] <= 1;
      stuckIsFree_memory[5] <= 1;
      stuckIsFree_memory[6] <= 1;
      stuckIsFree_memory[7] <= 1;
      stuckIsFree_memory[8] <= 1;
      stuckIsFree_memory[9] <= 1;
      stuckIsFree_memory[10] <= 1;
      stuckIsFree_memory[11] <= 1;
      stuckIsFree_memory[12] <= 1;
      stuckIsFree_memory[13] <= 1;
      stuckIsFree_memory[14] <= 1;
      stuckIsFree_memory[15] <= 1;
      stuckIsFree_memory[16] <= 1;
      stuckIsFree_memory[17] <= 1;
      stuckIsFree_memory[18] <= 1;
      stuckIsFree_memory[19] <= 1;
      stuckIsFree_memory[20] <= 1;
      stuckIsFree_memory[21] <= 1;
      stuckIsFree_memory[22] <= 1;
      stuckIsFree_memory[23] <= 1;
      stuckIsFree_memory[24] <= 1;
      stuckIsFree_memory[25] <= 1;
      stuckIsFree_memory[26] <= 1;
      stuckIsFree_memory[27] <= 1;
      stuckIsFree_memory[28] <= 1;
      stuckIsFree_memory[29] <= 1;
      stuckIsFree_memory[30] <= 1;
      stuckIsFree_memory[31] <= 1;
    end
    else if (processCurrent == 1) begin
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step)) begin
            stuckIsFree_memory[findAndInsert_stuckIsFree_11_index_171*1+0] <= findAndInsert_stuckIsFree_11_value_172;
            stuckIsFree_11_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [6-1:0] freeNext_memory[32*1];
  reg [6-1:0] freeNext_freeNext_9_result_0;
  integer freeNext_9_requestedAt;
  integer freeNext_9_finishedAt;
  integer freeNext_freeNext_9_returnCode;
  integer freeNext_10_requestedAt;
  integer freeNext_10_finishedAt;
  integer freeNext_freeNext_10_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_9_result_0 <= 0;
      freeNext_9_finishedAt <= -1;
      freeNext_freeNext_9_returnCode <= 0;
      freeNext_10_finishedAt <= -1;
      freeNext_freeNext_10_returnCode <= 0;
      freeNext_memory[0] <= 1;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 7;
      freeNext_memory[7] <= 8;
      freeNext_memory[8] <= 9;
      freeNext_memory[9] <= 10;
      freeNext_memory[10] <= 11;
      freeNext_memory[11] <= 12;
      freeNext_memory[12] <= 13;
      freeNext_memory[13] <= 14;
      freeNext_memory[14] <= 15;
      freeNext_memory[15] <= 16;
      freeNext_memory[16] <= 17;
      freeNext_memory[17] <= 18;
      freeNext_memory[18] <= 19;
      freeNext_memory[19] <= 20;
      freeNext_memory[20] <= 21;
      freeNext_memory[21] <= 22;
      freeNext_memory[22] <= 23;
      freeNext_memory[23] <= 24;
      freeNext_memory[24] <= 25;
      freeNext_memory[25] <= 26;
      freeNext_memory[26] <= 27;
      freeNext_memory[27] <= 28;
      freeNext_memory[28] <= 29;
      freeNext_memory[29] <= 30;
      freeNext_memory[30] <= 31;
      freeNext_memory[31] <= 0;
    end
    else if (processCurrent == 2) begin
      case(freeNext_pc)
        0: begin
          if ((freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step)) begin
            freeNext_freeNext_9_result_0 <= freeNext_memory[findAndInsert_freeNext_9_index_168*1+0];
            freeNext_9_finishedAt <= step;
          end
          else if ((freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step)) begin
            freeNext_memory[findAndInsert_freeNext_10_index_169*1+0] <= findAndInsert_freeNext_10_value_170;
            freeNext_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[32*1];
  reg [3-1:0] stuckSize_stuckSize_5_result_0;
  integer stuckSize_5_requestedAt;
  integer stuckSize_5_finishedAt;
  integer stuckSize_stuckSize_5_returnCode;
  integer stuckSize_6_requestedAt;
  integer stuckSize_6_finishedAt;
  integer stuckSize_stuckSize_6_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_5_result_0 <= 0;
      stuckSize_5_finishedAt <= -1;
      stuckSize_stuckSize_5_returnCode <= 0;
      stuckSize_6_finishedAt <= -1;
      stuckSize_stuckSize_6_returnCode <= 0;
      stuckSize_memory[0] <= 0;
      stuckSize_memory[1] <= 0;
      stuckSize_memory[2] <= 0;
      stuckSize_memory[3] <= 0;
      stuckSize_memory[4] <= 0;
      stuckSize_memory[5] <= 0;
      stuckSize_memory[6] <= 0;
      stuckSize_memory[7] <= 0;
      stuckSize_memory[8] <= 0;
      stuckSize_memory[9] <= 0;
      stuckSize_memory[10] <= 0;
      stuckSize_memory[11] <= 0;
      stuckSize_memory[12] <= 0;
      stuckSize_memory[13] <= 0;
      stuckSize_memory[14] <= 0;
      stuckSize_memory[15] <= 0;
      stuckSize_memory[16] <= 0;
      stuckSize_memory[17] <= 0;
      stuckSize_memory[18] <= 0;
      stuckSize_memory[19] <= 0;
      stuckSize_memory[20] <= 0;
      stuckSize_memory[21] <= 0;
      stuckSize_memory[22] <= 0;
      stuckSize_memory[23] <= 0;
      stuckSize_memory[24] <= 0;
      stuckSize_memory[25] <= 0;
      stuckSize_memory[26] <= 0;
      stuckSize_memory[27] <= 0;
      stuckSize_memory[28] <= 0;
      stuckSize_memory[29] <= 0;
      stuckSize_memory[30] <= 0;
      stuckSize_memory[31] <= 0;
    end
    else if (processCurrent == 3) begin
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step)) begin
            stuckSize_stuckSize_5_result_0 <= stuckSize_memory[findAndInsert_stuckSize_5_index_32*1+0];
            stuckSize_5_finishedAt <= step;
          end
          else if ((stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step)) begin
            stuckSize_memory[findAndInsert_stuckSize_6_index_33*1+0] <= findAndInsert_stuckSize_6_value_34;
            stuckSize_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys  process_stuckKeys_0004
  (* ram_style = "block" *)
  reg [8-1:0] stuckKeys_memory[32*4];
  reg [8-1:0] stuckKeys_stuckKeys_1_result_0;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_1;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_2;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_3;
  integer stuckKeys_1_requestedAt;
  integer stuckKeys_1_finishedAt;
  integer stuckKeys_stuckKeys_1_returnCode;
  integer stuckKeys_2_requestedAt;
  integer stuckKeys_2_finishedAt;
  integer stuckKeys_stuckKeys_2_returnCode;
  integer stuckKeys_pc;
  integer stuckKeys_stop;
  integer stuckKeys_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_pc <= 0;
      stuckKeys_stop <= 0;
      stuckKeys_returnCode <= 0;
      stuckKeys_stuckKeys_1_result_0 <= 0;
      stuckKeys_stuckKeys_1_result_1 <= 0;
      stuckKeys_stuckKeys_1_result_2 <= 0;
      stuckKeys_stuckKeys_1_result_3 <= 0;
      stuckKeys_1_finishedAt <= -1;
      stuckKeys_stuckKeys_1_returnCode <= 0;
      stuckKeys_2_finishedAt <= -1;
      stuckKeys_stuckKeys_2_returnCode <= 0;
      stuckKeys_memory[0] <= 0;
      stuckKeys_memory[1] <= 0;
      stuckKeys_memory[2] <= 0;
      stuckKeys_memory[3] <= 0;
      stuckKeys_memory[4] <= 0;
      stuckKeys_memory[5] <= 0;
      stuckKeys_memory[6] <= 0;
      stuckKeys_memory[7] <= 0;
      stuckKeys_memory[8] <= 0;
      stuckKeys_memory[9] <= 0;
      stuckKeys_memory[10] <= 0;
      stuckKeys_memory[11] <= 0;
      stuckKeys_memory[12] <= 0;
      stuckKeys_memory[13] <= 0;
      stuckKeys_memory[14] <= 0;
      stuckKeys_memory[15] <= 0;
      stuckKeys_memory[16] <= 0;
      stuckKeys_memory[17] <= 0;
      stuckKeys_memory[18] <= 0;
      stuckKeys_memory[19] <= 0;
      stuckKeys_memory[20] <= 0;
      stuckKeys_memory[21] <= 0;
      stuckKeys_memory[22] <= 0;
      stuckKeys_memory[23] <= 0;
      stuckKeys_memory[24] <= 0;
      stuckKeys_memory[25] <= 0;
      stuckKeys_memory[26] <= 0;
      stuckKeys_memory[27] <= 0;
      stuckKeys_memory[28] <= 0;
      stuckKeys_memory[29] <= 0;
      stuckKeys_memory[30] <= 0;
      stuckKeys_memory[31] <= 0;
      stuckKeys_memory[32] <= 0;
      stuckKeys_memory[33] <= 0;
      stuckKeys_memory[34] <= 0;
      stuckKeys_memory[35] <= 0;
      stuckKeys_memory[36] <= 0;
      stuckKeys_memory[37] <= 0;
      stuckKeys_memory[38] <= 0;
      stuckKeys_memory[39] <= 0;
      stuckKeys_memory[40] <= 0;
      stuckKeys_memory[41] <= 0;
      stuckKeys_memory[42] <= 0;
      stuckKeys_memory[43] <= 0;
      stuckKeys_memory[44] <= 0;
      stuckKeys_memory[45] <= 0;
      stuckKeys_memory[46] <= 0;
      stuckKeys_memory[47] <= 0;
      stuckKeys_memory[48] <= 0;
      stuckKeys_memory[49] <= 0;
      stuckKeys_memory[50] <= 0;
      stuckKeys_memory[51] <= 0;
      stuckKeys_memory[52] <= 0;
      stuckKeys_memory[53] <= 0;
      stuckKeys_memory[54] <= 0;
      stuckKeys_memory[55] <= 0;
      stuckKeys_memory[56] <= 0;
      stuckKeys_memory[57] <= 0;
      stuckKeys_memory[58] <= 0;
      stuckKeys_memory[59] <= 0;
      stuckKeys_memory[60] <= 0;
      stuckKeys_memory[61] <= 0;
      stuckKeys_memory[62] <= 0;
      stuckKeys_memory[63] <= 0;
      stuckKeys_memory[64] <= 0;
      stuckKeys_memory[65] <= 0;
      stuckKeys_memory[66] <= 0;
      stuckKeys_memory[67] <= 0;
      stuckKeys_memory[68] <= 0;
      stuckKeys_memory[69] <= 0;
      stuckKeys_memory[70] <= 0;
      stuckKeys_memory[71] <= 0;
      stuckKeys_memory[72] <= 0;
      stuckKeys_memory[73] <= 0;
      stuckKeys_memory[74] <= 0;
      stuckKeys_memory[75] <= 0;
      stuckKeys_memory[76] <= 0;
      stuckKeys_memory[77] <= 0;
      stuckKeys_memory[78] <= 0;
      stuckKeys_memory[79] <= 0;
      stuckKeys_memory[80] <= 0;
      stuckKeys_memory[81] <= 0;
      stuckKeys_memory[82] <= 0;
      stuckKeys_memory[83] <= 0;
      stuckKeys_memory[84] <= 0;
      stuckKeys_memory[85] <= 0;
      stuckKeys_memory[86] <= 0;
      stuckKeys_memory[87] <= 0;
      stuckKeys_memory[88] <= 0;
      stuckKeys_memory[89] <= 0;
      stuckKeys_memory[90] <= 0;
      stuckKeys_memory[91] <= 0;
      stuckKeys_memory[92] <= 0;
      stuckKeys_memory[93] <= 0;
      stuckKeys_memory[94] <= 0;
      stuckKeys_memory[95] <= 0;
      stuckKeys_memory[96] <= 0;
      stuckKeys_memory[97] <= 0;
      stuckKeys_memory[98] <= 0;
      stuckKeys_memory[99] <= 0;
      stuckKeys_memory[100] <= 0;
      stuckKeys_memory[101] <= 0;
      stuckKeys_memory[102] <= 0;
      stuckKeys_memory[103] <= 0;
      stuckKeys_memory[104] <= 0;
      stuckKeys_memory[105] <= 0;
      stuckKeys_memory[106] <= 0;
      stuckKeys_memory[107] <= 0;
      stuckKeys_memory[108] <= 0;
      stuckKeys_memory[109] <= 0;
      stuckKeys_memory[110] <= 0;
      stuckKeys_memory[111] <= 0;
      stuckKeys_memory[112] <= 0;
      stuckKeys_memory[113] <= 0;
      stuckKeys_memory[114] <= 0;
      stuckKeys_memory[115] <= 0;
      stuckKeys_memory[116] <= 0;
      stuckKeys_memory[117] <= 0;
      stuckKeys_memory[118] <= 0;
      stuckKeys_memory[119] <= 0;
      stuckKeys_memory[120] <= 0;
      stuckKeys_memory[121] <= 0;
      stuckKeys_memory[122] <= 0;
      stuckKeys_memory[123] <= 0;
      stuckKeys_memory[124] <= 0;
      stuckKeys_memory[125] <= 0;
      stuckKeys_memory[126] <= 0;
      stuckKeys_memory[127] <= 0;
    end
    else if (processCurrent == 4) begin
      case(stuckKeys_pc)
        0: begin
          if ((stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step)) begin
            stuckKeys_stuckKeys_1_result_0 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+0];
            stuckKeys_stuckKeys_1_result_1 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+1];
            stuckKeys_stuckKeys_1_result_2 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+2];
            stuckKeys_stuckKeys_1_result_3 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+3];
            stuckKeys_1_finishedAt <= step;
          end
          else if ((stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step)) begin
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+0] <= findAndInsert_stuckKeys_2_value_22;
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+1] <= findAndInsert_stuckKeys_2_value_23;
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+2] <= findAndInsert_stuckKeys_2_value_24;
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+3] <= findAndInsert_stuckKeys_2_value_25;
            stuckKeys_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_stop <= 1;
      endcase
    end
  end
  // Process: stuckData  process_stuckData_0005
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_memory[32*4];
  reg [8-1:0] stuckData_stuckData_3_result_0;
  reg [8-1:0] stuckData_stuckData_3_result_1;
  reg [8-1:0] stuckData_stuckData_3_result_2;
  reg [8-1:0] stuckData_stuckData_3_result_3;
  integer stuckData_3_requestedAt;
  integer stuckData_3_finishedAt;
  integer stuckData_stuckData_3_returnCode;
  integer stuckData_4_requestedAt;
  integer stuckData_4_finishedAt;
  integer stuckData_stuckData_4_returnCode;
  integer stuckData_pc;
  integer stuckData_stop;
  integer stuckData_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_pc <= 0;
      stuckData_stop <= 0;
      stuckData_returnCode <= 0;
      stuckData_stuckData_3_result_0 <= 0;
      stuckData_stuckData_3_result_1 <= 0;
      stuckData_stuckData_3_result_2 <= 0;
      stuckData_stuckData_3_result_3 <= 0;
      stuckData_3_finishedAt <= -1;
      stuckData_stuckData_3_returnCode <= 0;
      stuckData_4_finishedAt <= -1;
      stuckData_stuckData_4_returnCode <= 0;
      stuckData_memory[0] <= 0;
      stuckData_memory[1] <= 0;
      stuckData_memory[2] <= 0;
      stuckData_memory[3] <= 0;
      stuckData_memory[4] <= 0;
      stuckData_memory[5] <= 0;
      stuckData_memory[6] <= 0;
      stuckData_memory[7] <= 0;
      stuckData_memory[8] <= 0;
      stuckData_memory[9] <= 0;
      stuckData_memory[10] <= 0;
      stuckData_memory[11] <= 0;
      stuckData_memory[12] <= 0;
      stuckData_memory[13] <= 0;
      stuckData_memory[14] <= 0;
      stuckData_memory[15] <= 0;
      stuckData_memory[16] <= 0;
      stuckData_memory[17] <= 0;
      stuckData_memory[18] <= 0;
      stuckData_memory[19] <= 0;
      stuckData_memory[20] <= 0;
      stuckData_memory[21] <= 0;
      stuckData_memory[22] <= 0;
      stuckData_memory[23] <= 0;
      stuckData_memory[24] <= 0;
      stuckData_memory[25] <= 0;
      stuckData_memory[26] <= 0;
      stuckData_memory[27] <= 0;
      stuckData_memory[28] <= 0;
      stuckData_memory[29] <= 0;
      stuckData_memory[30] <= 0;
      stuckData_memory[31] <= 0;
      stuckData_memory[32] <= 0;
      stuckData_memory[33] <= 0;
      stuckData_memory[34] <= 0;
      stuckData_memory[35] <= 0;
      stuckData_memory[36] <= 0;
      stuckData_memory[37] <= 0;
      stuckData_memory[38] <= 0;
      stuckData_memory[39] <= 0;
      stuckData_memory[40] <= 0;
      stuckData_memory[41] <= 0;
      stuckData_memory[42] <= 0;
      stuckData_memory[43] <= 0;
      stuckData_memory[44] <= 0;
      stuckData_memory[45] <= 0;
      stuckData_memory[46] <= 0;
      stuckData_memory[47] <= 0;
      stuckData_memory[48] <= 0;
      stuckData_memory[49] <= 0;
      stuckData_memory[50] <= 0;
      stuckData_memory[51] <= 0;
      stuckData_memory[52] <= 0;
      stuckData_memory[53] <= 0;
      stuckData_memory[54] <= 0;
      stuckData_memory[55] <= 0;
      stuckData_memory[56] <= 0;
      stuckData_memory[57] <= 0;
      stuckData_memory[58] <= 0;
      stuckData_memory[59] <= 0;
      stuckData_memory[60] <= 0;
      stuckData_memory[61] <= 0;
      stuckData_memory[62] <= 0;
      stuckData_memory[63] <= 0;
      stuckData_memory[64] <= 0;
      stuckData_memory[65] <= 0;
      stuckData_memory[66] <= 0;
      stuckData_memory[67] <= 0;
      stuckData_memory[68] <= 0;
      stuckData_memory[69] <= 0;
      stuckData_memory[70] <= 0;
      stuckData_memory[71] <= 0;
      stuckData_memory[72] <= 0;
      stuckData_memory[73] <= 0;
      stuckData_memory[74] <= 0;
      stuckData_memory[75] <= 0;
      stuckData_memory[76] <= 0;
      stuckData_memory[77] <= 0;
      stuckData_memory[78] <= 0;
      stuckData_memory[79] <= 0;
      stuckData_memory[80] <= 0;
      stuckData_memory[81] <= 0;
      stuckData_memory[82] <= 0;
      stuckData_memory[83] <= 0;
      stuckData_memory[84] <= 0;
      stuckData_memory[85] <= 0;
      stuckData_memory[86] <= 0;
      stuckData_memory[87] <= 0;
      stuckData_memory[88] <= 0;
      stuckData_memory[89] <= 0;
      stuckData_memory[90] <= 0;
      stuckData_memory[91] <= 0;
      stuckData_memory[92] <= 0;
      stuckData_memory[93] <= 0;
      stuckData_memory[94] <= 0;
      stuckData_memory[95] <= 0;
      stuckData_memory[96] <= 0;
      stuckData_memory[97] <= 0;
      stuckData_memory[98] <= 0;
      stuckData_memory[99] <= 0;
      stuckData_memory[100] <= 0;
      stuckData_memory[101] <= 0;
      stuckData_memory[102] <= 0;
      stuckData_memory[103] <= 0;
      stuckData_memory[104] <= 0;
      stuckData_memory[105] <= 0;
      stuckData_memory[106] <= 0;
      stuckData_memory[107] <= 0;
      stuckData_memory[108] <= 0;
      stuckData_memory[109] <= 0;
      stuckData_memory[110] <= 0;
      stuckData_memory[111] <= 0;
      stuckData_memory[112] <= 0;
      stuckData_memory[113] <= 0;
      stuckData_memory[114] <= 0;
      stuckData_memory[115] <= 0;
      stuckData_memory[116] <= 0;
      stuckData_memory[117] <= 0;
      stuckData_memory[118] <= 0;
      stuckData_memory[119] <= 0;
      stuckData_memory[120] <= 0;
      stuckData_memory[121] <= 0;
      stuckData_memory[122] <= 0;
      stuckData_memory[123] <= 0;
      stuckData_memory[124] <= 0;
      stuckData_memory[125] <= 0;
      stuckData_memory[126] <= 0;
      stuckData_memory[127] <= 0;
    end
    else if (processCurrent == 5) begin
      case(stuckData_pc)
        0: begin
          if ((stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step)) begin
            stuckData_stuckData_3_result_0 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+0];
            stuckData_stuckData_3_result_1 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+1];
            stuckData_stuckData_3_result_2 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+2];
            stuckData_stuckData_3_result_3 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+3];
            stuckData_3_finishedAt <= step;
          end
          else if ((stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step)) begin
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+0] <= findAndInsert_stuckData_4_value_28;
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+1] <= findAndInsert_stuckData_4_value_29;
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+2] <= findAndInsert_stuckData_4_value_30;
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+3] <= findAndInsert_stuckData_4_value_31;
            stuckData_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_stop <= 1;
      endcase
    end
  end
  // Process: findAndInsert  process_findAndInsert_0006
  reg [6-1:0] findAndInsert_index_0;
  reg [3-1:0] findAndInsert_size_1;
  reg [1-1:0] findAndInsert_isLeaf_2;
  reg [6-1:0] findAndInsert_nextFree_3;
  reg [8-1:0] findAndInsert_Key_0_4;
  reg [1-1:0] findAndInsert_KeyCompares_0_5;
  reg [3-1:0] findAndInsert_KeyCollapse_0_6;
  reg [8-1:0] findAndInsert_Data_0_7;
  reg [8-1:0] findAndInsert_Key_1_8;
  reg [1-1:0] findAndInsert_KeyCompares_1_9;
  reg [3-1:0] findAndInsert_KeyCollapse_1_10;
  reg [8-1:0] findAndInsert_Data_1_11;
  reg [8-1:0] findAndInsert_Key_2_12;
  reg [1-1:0] findAndInsert_KeyCompares_2_13;
  reg [3-1:0] findAndInsert_KeyCollapse_2_14;
  reg [8-1:0] findAndInsert_Data_2_15;
  reg [8-1:0] findAndInsert_Key_3_16;
  reg [1-1:0] findAndInsert_KeyCompares_3_17;
  reg [3-1:0] findAndInsert_KeyCollapse_3_18;
  reg [8-1:0] findAndInsert_Data_3_19;
  reg [5-1:0] findAndInsert_stuckKeys_1_index_20;
  reg [5-1:0] findAndInsert_stuckKeys_2_index_21;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_22;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_23;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_24;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_25;
  reg [5-1:0] findAndInsert_stuckData_3_index_26;
  reg [5-1:0] findAndInsert_stuckData_4_index_27;
  reg [8-1:0] findAndInsert_stuckData_4_value_28;
  reg [8-1:0] findAndInsert_stuckData_4_value_29;
  reg [8-1:0] findAndInsert_stuckData_4_value_30;
  reg [8-1:0] findAndInsert_stuckData_4_value_31;
  reg [5-1:0] findAndInsert_stuckSize_5_index_32;
  reg [5-1:0] findAndInsert_stuckSize_6_index_33;
  reg [3-1:0] findAndInsert_stuckSize_6_value_34;
  reg [5-1:0] findAndInsert_stuckIsLeaf_7_index_35;
  reg [5-1:0] findAndInsert_stuckIsLeaf_8_index_36;
  reg [1-1:0] findAndInsert_stuckIsLeaf_8_value_37;
  reg [1-1:0] findAndInsert_Found_38;
  reg [8-1:0] findAndInsert_Key_39;
  reg [8-1:0] findAndInsert_FoundKey_40;
  reg [8-1:0] findAndInsert_Data_41;
  reg [6-1:0] findAndInsert_BtreeIndex_42;
  reg [3-1:0] findAndInsert_StuckIndex_43;
  reg [1-1:0] findAndInsert_MergeSuccess_44;
  reg [8-1:0] findAndInsert_k_45;
  reg [8-1:0] findAndInsert_d_46;
  reg [6-1:0] findAndInsert_i_47;
  reg [3-1:0] findAndInsert_j_48;
  reg [6-1:0] findAndInsert_index_49;
  reg [3-1:0] findAndInsert_size_50;
  reg [1-1:0] findAndInsert_isLeaf_51;
  reg [6-1:0] findAndInsert_nextFree_52;
  reg [8-1:0] findAndInsert_Key_0_53;
  reg [1-1:0] findAndInsert_KeyCompares_0_54;
  reg [3-1:0] findAndInsert_KeyCollapse_0_55;
  reg [8-1:0] findAndInsert_Data_0_56;
  reg [8-1:0] findAndInsert_Key_1_57;
  reg [1-1:0] findAndInsert_KeyCompares_1_58;
  reg [3-1:0] findAndInsert_KeyCollapse_1_59;
  reg [8-1:0] findAndInsert_Data_1_60;
  reg [8-1:0] findAndInsert_Key_2_61;
  reg [1-1:0] findAndInsert_KeyCompares_2_62;
  reg [3-1:0] findAndInsert_KeyCollapse_2_63;
  reg [8-1:0] findAndInsert_Data_2_64;
  reg [8-1:0] findAndInsert_Key_3_65;
  reg [1-1:0] findAndInsert_KeyCompares_3_66;
  reg [3-1:0] findAndInsert_KeyCollapse_3_67;
  reg [8-1:0] findAndInsert_Data_3_68;
  reg [1-1:0] findAndInsert_Found_69;
  reg [8-1:0] findAndInsert_Key_70;
  reg [8-1:0] findAndInsert_FoundKey_71;
  reg [8-1:0] findAndInsert_Data_72;
  reg [6-1:0] findAndInsert_BtreeIndex_73;
  reg [3-1:0] findAndInsert_StuckIndex_74;
  reg [1-1:0] findAndInsert_MergeSuccess_75;
  reg [3-1:0] findAndInsert_i_76;
  reg [1-1:0] findAndInsert_notFull_77;
  reg [3-1:0] findAndInsert_i_78;
  reg [1-1:0] findAndInsert_notFull_79;
  reg [3-1:0] findAndInsert_i_80;
  reg [1-1:0] findAndInsert_notFull_81;
  reg [3-1:0] findAndInsert_i_82;
  reg [1-1:0] findAndInsert_notFull_83;
  reg [6-1:0] findAndInsert_index_84;
  reg [3-1:0] findAndInsert_size_85;
  reg [1-1:0] findAndInsert_isLeaf_86;
  reg [6-1:0] findAndInsert_nextFree_87;
  reg [8-1:0] findAndInsert_Key_0_88;
  reg [1-1:0] findAndInsert_KeyCompares_0_89;
  reg [3-1:0] findAndInsert_KeyCollapse_0_90;
  reg [8-1:0] findAndInsert_Data_0_91;
  reg [8-1:0] findAndInsert_Key_1_92;
  reg [1-1:0] findAndInsert_KeyCompares_1_93;
  reg [3-1:0] findAndInsert_KeyCollapse_1_94;
  reg [8-1:0] findAndInsert_Data_1_95;
  reg [8-1:0] findAndInsert_Key_2_96;
  reg [1-1:0] findAndInsert_KeyCompares_2_97;
  reg [3-1:0] findAndInsert_KeyCollapse_2_98;
  reg [8-1:0] findAndInsert_Data_2_99;
  reg [8-1:0] findAndInsert_Key_3_100;
  reg [1-1:0] findAndInsert_KeyCompares_3_101;
  reg [3-1:0] findAndInsert_KeyCollapse_3_102;
  reg [8-1:0] findAndInsert_Data_3_103;
  reg [1-1:0] findAndInsert_Found_104;
  reg [8-1:0] findAndInsert_Key_105;
  reg [8-1:0] findAndInsert_FoundKey_106;
  reg [8-1:0] findAndInsert_Data_107;
  reg [6-1:0] findAndInsert_BtreeIndex_108;
  reg [3-1:0] findAndInsert_StuckIndex_109;
  reg [1-1:0] findAndInsert_MergeSuccess_110;
  reg [6-1:0] findAndInsert_index_111;
  reg [3-1:0] findAndInsert_size_112;
  reg [1-1:0] findAndInsert_isLeaf_113;
  reg [6-1:0] findAndInsert_nextFree_114;
  reg [8-1:0] findAndInsert_Key_0_115;
  reg [1-1:0] findAndInsert_KeyCompares_0_116;
  reg [3-1:0] findAndInsert_KeyCollapse_0_117;
  reg [8-1:0] findAndInsert_Data_0_118;
  reg [8-1:0] findAndInsert_Key_1_119;
  reg [1-1:0] findAndInsert_KeyCompares_1_120;
  reg [3-1:0] findAndInsert_KeyCollapse_1_121;
  reg [8-1:0] findAndInsert_Data_1_122;
  reg [8-1:0] findAndInsert_Key_2_123;
  reg [1-1:0] findAndInsert_KeyCompares_2_124;
  reg [3-1:0] findAndInsert_KeyCollapse_2_125;
  reg [8-1:0] findAndInsert_Data_2_126;
  reg [8-1:0] findAndInsert_Key_3_127;
  reg [1-1:0] findAndInsert_KeyCompares_3_128;
  reg [3-1:0] findAndInsert_KeyCollapse_3_129;
  reg [8-1:0] findAndInsert_Data_3_130;
  reg [1-1:0] findAndInsert_Found_131;
  reg [8-1:0] findAndInsert_Key_132;
  reg [8-1:0] findAndInsert_FoundKey_133;
  reg [8-1:0] findAndInsert_Data_134;
  reg [6-1:0] findAndInsert_BtreeIndex_135;
  reg [3-1:0] findAndInsert_StuckIndex_136;
  reg [1-1:0] findAndInsert_MergeSuccess_137;
  reg [6-1:0] findAndInsert_index_138;
  reg [3-1:0] findAndInsert_size_139;
  reg [1-1:0] findAndInsert_isLeaf_140;
  reg [6-1:0] findAndInsert_nextFree_141;
  reg [8-1:0] findAndInsert_Key_0_142;
  reg [1-1:0] findAndInsert_KeyCompares_0_143;
  reg [3-1:0] findAndInsert_KeyCollapse_0_144;
  reg [8-1:0] findAndInsert_Data_0_145;
  reg [8-1:0] findAndInsert_Key_1_146;
  reg [1-1:0] findAndInsert_KeyCompares_1_147;
  reg [3-1:0] findAndInsert_KeyCollapse_1_148;
  reg [8-1:0] findAndInsert_Data_1_149;
  reg [8-1:0] findAndInsert_Key_2_150;
  reg [1-1:0] findAndInsert_KeyCompares_2_151;
  reg [3-1:0] findAndInsert_KeyCollapse_2_152;
  reg [8-1:0] findAndInsert_Data_2_153;
  reg [8-1:0] findAndInsert_Key_3_154;
  reg [1-1:0] findAndInsert_KeyCompares_3_155;
  reg [3-1:0] findAndInsert_KeyCollapse_3_156;
  reg [8-1:0] findAndInsert_Data_3_157;
  reg [1-1:0] findAndInsert_Found_158;
  reg [8-1:0] findAndInsert_Key_159;
  reg [8-1:0] findAndInsert_FoundKey_160;
  reg [8-1:0] findAndInsert_Data_161;
  reg [6-1:0] findAndInsert_BtreeIndex_162;
  reg [3-1:0] findAndInsert_StuckIndex_163;
  reg [1-1:0] findAndInsert_MergeSuccess_164;
  reg [6-1:0] findAndInsert_indexLeft_165;
  reg [6-1:0] findAndInsert_indexRight_166;
  reg [8-1:0] findAndInsert_midKey_167;
  reg [5-1:0] findAndInsert_freeNext_9_index_168;
  reg [5-1:0] findAndInsert_freeNext_10_index_169;
  reg [6-1:0] findAndInsert_freeNext_10_value_170;
  reg [5-1:0] findAndInsert_stuckIsFree_11_index_171;
  reg [1-1:0] findAndInsert_stuckIsFree_11_value_172;
  reg [6-1:0] findAndInsert_root_173;
  reg [6-1:0] findAndInsert_next_174;
  reg [1-1:0] findAndInsert_isLeaf_175;
  reg [1-1:0] findAndInsert_isFree_176;
  reg [6-1:0] findAndInsert_root_177;
  reg [6-1:0] findAndInsert_next_178;
  reg [1-1:0] findAndInsert_isLeaf_179;
  reg [1-1:0] findAndInsert_isFree_180;
  reg [3-1:0] findAndInsert_i_181;
  reg [1-1:0] findAndInsert_notFull_182;
  reg [3-1:0] findAndInsert_i_183;
  reg [1-1:0] findAndInsert_notFull_184;
  reg [6-1:0] findAndInsert_index_185;
  reg [3-1:0] findAndInsert_size_186;
  reg [1-1:0] findAndInsert_isLeaf_187;
  reg [6-1:0] findAndInsert_nextFree_188;
  reg [8-1:0] findAndInsert_Key_0_189;
  reg [1-1:0] findAndInsert_KeyCompares_0_190;
  reg [3-1:0] findAndInsert_KeyCollapse_0_191;
  reg [8-1:0] findAndInsert_Data_0_192;
  reg [8-1:0] findAndInsert_Key_1_193;
  reg [1-1:0] findAndInsert_KeyCompares_1_194;
  reg [3-1:0] findAndInsert_KeyCollapse_1_195;
  reg [8-1:0] findAndInsert_Data_1_196;
  reg [8-1:0] findAndInsert_Key_2_197;
  reg [1-1:0] findAndInsert_KeyCompares_2_198;
  reg [3-1:0] findAndInsert_KeyCollapse_2_199;
  reg [8-1:0] findAndInsert_Data_2_200;
  reg [8-1:0] findAndInsert_Key_3_201;
  reg [1-1:0] findAndInsert_KeyCompares_3_202;
  reg [3-1:0] findAndInsert_KeyCollapse_3_203;
  reg [8-1:0] findAndInsert_Data_3_204;
  reg [1-1:0] findAndInsert_Found_205;
  reg [8-1:0] findAndInsert_Key_206;
  reg [8-1:0] findAndInsert_FoundKey_207;
  reg [8-1:0] findAndInsert_Data_208;
  reg [6-1:0] findAndInsert_BtreeIndex_209;
  reg [3-1:0] findAndInsert_StuckIndex_210;
  reg [1-1:0] findAndInsert_MergeSuccess_211;
  reg [6-1:0] findAndInsert_index_212;
  reg [3-1:0] findAndInsert_size_213;
  reg [1-1:0] findAndInsert_isLeaf_214;
  reg [6-1:0] findAndInsert_nextFree_215;
  reg [8-1:0] findAndInsert_Key_0_216;
  reg [1-1:0] findAndInsert_KeyCompares_0_217;
  reg [3-1:0] findAndInsert_KeyCollapse_0_218;
  reg [8-1:0] findAndInsert_Data_0_219;
  reg [8-1:0] findAndInsert_Key_1_220;
  reg [1-1:0] findAndInsert_KeyCompares_1_221;
  reg [3-1:0] findAndInsert_KeyCollapse_1_222;
  reg [8-1:0] findAndInsert_Data_1_223;
  reg [8-1:0] findAndInsert_Key_2_224;
  reg [1-1:0] findAndInsert_KeyCompares_2_225;
  reg [3-1:0] findAndInsert_KeyCollapse_2_226;
  reg [8-1:0] findAndInsert_Data_2_227;
  reg [8-1:0] findAndInsert_Key_3_228;
  reg [1-1:0] findAndInsert_KeyCompares_3_229;
  reg [3-1:0] findAndInsert_KeyCollapse_3_230;
  reg [8-1:0] findAndInsert_Data_3_231;
  reg [1-1:0] findAndInsert_Found_232;
  reg [8-1:0] findAndInsert_Key_233;
  reg [8-1:0] findAndInsert_FoundKey_234;
  reg [8-1:0] findAndInsert_Data_235;
  reg [6-1:0] findAndInsert_BtreeIndex_236;
  reg [3-1:0] findAndInsert_StuckIndex_237;
  reg [1-1:0] findAndInsert_MergeSuccess_238;
  reg [6-1:0] findAndInsert_index_239;
  reg [3-1:0] findAndInsert_size_240;
  reg [1-1:0] findAndInsert_isLeaf_241;
  reg [6-1:0] findAndInsert_nextFree_242;
  reg [8-1:0] findAndInsert_Key_0_243;
  reg [1-1:0] findAndInsert_KeyCompares_0_244;
  reg [3-1:0] findAndInsert_KeyCollapse_0_245;
  reg [8-1:0] findAndInsert_Data_0_246;
  reg [8-1:0] findAndInsert_Key_1_247;
  reg [1-1:0] findAndInsert_KeyCompares_1_248;
  reg [3-1:0] findAndInsert_KeyCollapse_1_249;
  reg [8-1:0] findAndInsert_Data_1_250;
  reg [8-1:0] findAndInsert_Key_2_251;
  reg [1-1:0] findAndInsert_KeyCompares_2_252;
  reg [3-1:0] findAndInsert_KeyCollapse_2_253;
  reg [8-1:0] findAndInsert_Data_2_254;
  reg [8-1:0] findAndInsert_Key_3_255;
  reg [1-1:0] findAndInsert_KeyCompares_3_256;
  reg [3-1:0] findAndInsert_KeyCollapse_3_257;
  reg [8-1:0] findAndInsert_Data_3_258;
  reg [1-1:0] findAndInsert_Found_259;
  reg [8-1:0] findAndInsert_Key_260;
  reg [8-1:0] findAndInsert_FoundKey_261;
  reg [8-1:0] findAndInsert_Data_262;
  reg [6-1:0] findAndInsert_BtreeIndex_263;
  reg [3-1:0] findAndInsert_StuckIndex_264;
  reg [1-1:0] findAndInsert_MergeSuccess_265;
  reg [6-1:0] findAndInsert_childIndex_266;
  reg [6-1:0] findAndInsert_leftIndex_267;
  reg [8-1:0] findAndInsert_midKey_268;
  reg [6-1:0] findAndInsert_root_269;
  reg [6-1:0] findAndInsert_next_270;
  reg [1-1:0] findAndInsert_isLeaf_271;
  reg [1-1:0] findAndInsert_isFree_272;
  reg [6-1:0] findAndInsert_index_273;
  reg [3-1:0] findAndInsert_size_274;
  reg [1-1:0] findAndInsert_isLeaf_275;
  reg [6-1:0] findAndInsert_nextFree_276;
  reg [8-1:0] findAndInsert_Key_0_277;
  reg [1-1:0] findAndInsert_KeyCompares_0_278;
  reg [3-1:0] findAndInsert_KeyCollapse_0_279;
  reg [8-1:0] findAndInsert_Data_0_280;
  reg [8-1:0] findAndInsert_Key_1_281;
  reg [1-1:0] findAndInsert_KeyCompares_1_282;
  reg [3-1:0] findAndInsert_KeyCollapse_1_283;
  reg [8-1:0] findAndInsert_Data_1_284;
  reg [8-1:0] findAndInsert_Key_2_285;
  reg [1-1:0] findAndInsert_KeyCompares_2_286;
  reg [3-1:0] findAndInsert_KeyCollapse_2_287;
  reg [8-1:0] findAndInsert_Data_2_288;
  reg [8-1:0] findAndInsert_Key_3_289;
  reg [1-1:0] findAndInsert_KeyCompares_3_290;
  reg [3-1:0] findAndInsert_KeyCollapse_3_291;
  reg [8-1:0] findAndInsert_Data_3_292;
  reg [1-1:0] findAndInsert_Found_293;
  reg [8-1:0] findAndInsert_Key_294;
  reg [8-1:0] findAndInsert_FoundKey_295;
  reg [8-1:0] findAndInsert_Data_296;
  reg [6-1:0] findAndInsert_BtreeIndex_297;
  reg [3-1:0] findAndInsert_StuckIndex_298;
  reg [1-1:0] findAndInsert_MergeSuccess_299;
  reg [6-1:0] findAndInsert_index_300;
  reg [3-1:0] findAndInsert_size_301;
  reg [1-1:0] findAndInsert_isLeaf_302;
  reg [6-1:0] findAndInsert_nextFree_303;
  reg [8-1:0] findAndInsert_Key_0_304;
  reg [1-1:0] findAndInsert_KeyCompares_0_305;
  reg [3-1:0] findAndInsert_KeyCollapse_0_306;
  reg [8-1:0] findAndInsert_Data_0_307;
  reg [8-1:0] findAndInsert_Key_1_308;
  reg [1-1:0] findAndInsert_KeyCompares_1_309;
  reg [3-1:0] findAndInsert_KeyCollapse_1_310;
  reg [8-1:0] findAndInsert_Data_1_311;
  reg [8-1:0] findAndInsert_Key_2_312;
  reg [1-1:0] findAndInsert_KeyCompares_2_313;
  reg [3-1:0] findAndInsert_KeyCollapse_2_314;
  reg [8-1:0] findAndInsert_Data_2_315;
  reg [8-1:0] findAndInsert_Key_3_316;
  reg [1-1:0] findAndInsert_KeyCompares_3_317;
  reg [3-1:0] findAndInsert_KeyCollapse_3_318;
  reg [8-1:0] findAndInsert_Data_3_319;
  reg [1-1:0] findAndInsert_Found_320;
  reg [8-1:0] findAndInsert_Key_321;
  reg [8-1:0] findAndInsert_FoundKey_322;
  reg [8-1:0] findAndInsert_Data_323;
  reg [6-1:0] findAndInsert_BtreeIndex_324;
  reg [3-1:0] findAndInsert_StuckIndex_325;
  reg [1-1:0] findAndInsert_MergeSuccess_326;
  reg [8-1:0] findAndInsert_childKey_327;
  reg [6-1:0] findAndInsert_childData_328;
  reg [6-1:0] findAndInsert_indexLeft_329;
  reg [6-1:0] findAndInsert_indexRight_330;
  reg [8-1:0] findAndInsert_midKey_331;
  reg [1-1:0] findAndInsert_success_332;
  reg [1-1:0] findAndInsert_test_333;
  reg [6-1:0] findAndInsert_next_334;
  reg [6-1:0] findAndInsert_root_335;
  reg [1-1:0] findAndInsert_isFree_336;
  integer findAndInsert_pc;
  integer findAndInsert_stop;
  integer findAndInsert_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      findAndInsert_pc <= 0;
      findAndInsert_stop <= 0;
      findAndInsert_returnCode <= 0;
      findAndInsert_index_0 <= 0;
      findAndInsert_size_1 <= 0;
      findAndInsert_isLeaf_2 <= 0;
      findAndInsert_nextFree_3 <= 0;
      findAndInsert_Key_0_4 <= 0;
      findAndInsert_KeyCompares_0_5 <= 0;
      findAndInsert_KeyCollapse_0_6 <= 0;
      findAndInsert_Data_0_7 <= 0;
      findAndInsert_Key_1_8 <= 0;
      findAndInsert_KeyCompares_1_9 <= 0;
      findAndInsert_KeyCollapse_1_10 <= 0;
      findAndInsert_Data_1_11 <= 0;
      findAndInsert_Key_2_12 <= 0;
      findAndInsert_KeyCompares_2_13 <= 0;
      findAndInsert_KeyCollapse_2_14 <= 0;
      findAndInsert_Data_2_15 <= 0;
      findAndInsert_Key_3_16 <= 0;
      findAndInsert_KeyCompares_3_17 <= 0;
      findAndInsert_KeyCollapse_3_18 <= 0;
      findAndInsert_Data_3_19 <= 0;
      findAndInsert_stuckKeys_1_index_20 <= 0;
      findAndInsert_stuckKeys_2_index_21 <= 0;
      findAndInsert_stuckKeys_2_value_22 <= 0;
      findAndInsert_stuckKeys_2_value_23 <= 0;
      findAndInsert_stuckKeys_2_value_24 <= 0;
      findAndInsert_stuckKeys_2_value_25 <= 0;
      findAndInsert_stuckData_3_index_26 <= 0;
      findAndInsert_stuckData_4_index_27 <= 0;
      findAndInsert_stuckData_4_value_28 <= 0;
      findAndInsert_stuckData_4_value_29 <= 0;
      findAndInsert_stuckData_4_value_30 <= 0;
      findAndInsert_stuckData_4_value_31 <= 0;
      findAndInsert_stuckSize_5_index_32 <= 0;
      findAndInsert_stuckSize_6_index_33 <= 0;
      findAndInsert_stuckSize_6_value_34 <= 0;
      findAndInsert_stuckIsLeaf_7_index_35 <= 0;
      findAndInsert_stuckIsLeaf_8_index_36 <= 0;
      findAndInsert_stuckIsLeaf_8_value_37 <= 0;
      findAndInsert_Found_38 <= 0;
      findAndInsert_Key_39 <= 0;
      findAndInsert_FoundKey_40 <= 0;
      findAndInsert_Data_41 <= 0;
      findAndInsert_BtreeIndex_42 <= 0;
      findAndInsert_StuckIndex_43 <= 0;
      findAndInsert_MergeSuccess_44 <= 0;
      findAndInsert_k_45 <= 0;
      findAndInsert_d_46 <= 0;
      findAndInsert_i_47 <= 0;
      findAndInsert_j_48 <= 0;
      findAndInsert_index_49 <= 0;
      findAndInsert_size_50 <= 0;
      findAndInsert_isLeaf_51 <= 0;
      findAndInsert_nextFree_52 <= 0;
      findAndInsert_Key_0_53 <= 0;
      findAndInsert_KeyCompares_0_54 <= 0;
      findAndInsert_KeyCollapse_0_55 <= 0;
      findAndInsert_Data_0_56 <= 0;
      findAndInsert_Key_1_57 <= 0;
      findAndInsert_KeyCompares_1_58 <= 0;
      findAndInsert_KeyCollapse_1_59 <= 0;
      findAndInsert_Data_1_60 <= 0;
      findAndInsert_Key_2_61 <= 0;
      findAndInsert_KeyCompares_2_62 <= 0;
      findAndInsert_KeyCollapse_2_63 <= 0;
      findAndInsert_Data_2_64 <= 0;
      findAndInsert_Key_3_65 <= 0;
      findAndInsert_KeyCompares_3_66 <= 0;
      findAndInsert_KeyCollapse_3_67 <= 0;
      findAndInsert_Data_3_68 <= 0;
      findAndInsert_Found_69 <= 0;
      findAndInsert_Key_70 <= 0;
      findAndInsert_FoundKey_71 <= 0;
      findAndInsert_Data_72 <= 0;
      findAndInsert_BtreeIndex_73 <= 0;
      findAndInsert_StuckIndex_74 <= 0;
      findAndInsert_MergeSuccess_75 <= 0;
      findAndInsert_i_76 <= 0;
      findAndInsert_notFull_77 <= 0;
      findAndInsert_i_78 <= 0;
      findAndInsert_notFull_79 <= 0;
      findAndInsert_i_80 <= 0;
      findAndInsert_notFull_81 <= 0;
      findAndInsert_i_82 <= 0;
      findAndInsert_notFull_83 <= 0;
      findAndInsert_index_84 <= 0;
      findAndInsert_size_85 <= 0;
      findAndInsert_isLeaf_86 <= 0;
      findAndInsert_nextFree_87 <= 0;
      findAndInsert_Key_0_88 <= 0;
      findAndInsert_KeyCompares_0_89 <= 0;
      findAndInsert_KeyCollapse_0_90 <= 0;
      findAndInsert_Data_0_91 <= 0;
      findAndInsert_Key_1_92 <= 0;
      findAndInsert_KeyCompares_1_93 <= 0;
      findAndInsert_KeyCollapse_1_94 <= 0;
      findAndInsert_Data_1_95 <= 0;
      findAndInsert_Key_2_96 <= 0;
      findAndInsert_KeyCompares_2_97 <= 0;
      findAndInsert_KeyCollapse_2_98 <= 0;
      findAndInsert_Data_2_99 <= 0;
      findAndInsert_Key_3_100 <= 0;
      findAndInsert_KeyCompares_3_101 <= 0;
      findAndInsert_KeyCollapse_3_102 <= 0;
      findAndInsert_Data_3_103 <= 0;
      findAndInsert_Found_104 <= 0;
      findAndInsert_Key_105 <= 0;
      findAndInsert_FoundKey_106 <= 0;
      findAndInsert_Data_107 <= 0;
      findAndInsert_BtreeIndex_108 <= 0;
      findAndInsert_StuckIndex_109 <= 0;
      findAndInsert_MergeSuccess_110 <= 0;
      findAndInsert_index_111 <= 0;
      findAndInsert_size_112 <= 0;
      findAndInsert_isLeaf_113 <= 0;
      findAndInsert_nextFree_114 <= 0;
      findAndInsert_Key_0_115 <= 0;
      findAndInsert_KeyCompares_0_116 <= 0;
      findAndInsert_KeyCollapse_0_117 <= 0;
      findAndInsert_Data_0_118 <= 0;
      findAndInsert_Key_1_119 <= 0;
      findAndInsert_KeyCompares_1_120 <= 0;
      findAndInsert_KeyCollapse_1_121 <= 0;
      findAndInsert_Data_1_122 <= 0;
      findAndInsert_Key_2_123 <= 0;
      findAndInsert_KeyCompares_2_124 <= 0;
      findAndInsert_KeyCollapse_2_125 <= 0;
      findAndInsert_Data_2_126 <= 0;
      findAndInsert_Key_3_127 <= 0;
      findAndInsert_KeyCompares_3_128 <= 0;
      findAndInsert_KeyCollapse_3_129 <= 0;
      findAndInsert_Data_3_130 <= 0;
      findAndInsert_Found_131 <= 0;
      findAndInsert_Key_132 <= 0;
      findAndInsert_FoundKey_133 <= 0;
      findAndInsert_Data_134 <= 0;
      findAndInsert_BtreeIndex_135 <= 0;
      findAndInsert_StuckIndex_136 <= 0;
      findAndInsert_MergeSuccess_137 <= 0;
      findAndInsert_index_138 <= 0;
      findAndInsert_size_139 <= 0;
      findAndInsert_isLeaf_140 <= 0;
      findAndInsert_nextFree_141 <= 0;
      findAndInsert_Key_0_142 <= 0;
      findAndInsert_KeyCompares_0_143 <= 0;
      findAndInsert_KeyCollapse_0_144 <= 0;
      findAndInsert_Data_0_145 <= 0;
      findAndInsert_Key_1_146 <= 0;
      findAndInsert_KeyCompares_1_147 <= 0;
      findAndInsert_KeyCollapse_1_148 <= 0;
      findAndInsert_Data_1_149 <= 0;
      findAndInsert_Key_2_150 <= 0;
      findAndInsert_KeyCompares_2_151 <= 0;
      findAndInsert_KeyCollapse_2_152 <= 0;
      findAndInsert_Data_2_153 <= 0;
      findAndInsert_Key_3_154 <= 0;
      findAndInsert_KeyCompares_3_155 <= 0;
      findAndInsert_KeyCollapse_3_156 <= 0;
      findAndInsert_Data_3_157 <= 0;
      findAndInsert_Found_158 <= 0;
      findAndInsert_Key_159 <= 0;
      findAndInsert_FoundKey_160 <= 0;
      findAndInsert_Data_161 <= 0;
      findAndInsert_BtreeIndex_162 <= 0;
      findAndInsert_StuckIndex_163 <= 0;
      findAndInsert_MergeSuccess_164 <= 0;
      findAndInsert_indexLeft_165 <= 0;
      findAndInsert_indexRight_166 <= 0;
      findAndInsert_midKey_167 <= 0;
      findAndInsert_freeNext_9_index_168 <= 0;
      findAndInsert_freeNext_10_index_169 <= 0;
      findAndInsert_freeNext_10_value_170 <= 0;
      findAndInsert_stuckIsFree_11_index_171 <= 0;
      findAndInsert_stuckIsFree_11_value_172 <= 0;
      findAndInsert_root_173 <= 0;
      findAndInsert_next_174 <= 0;
      findAndInsert_isLeaf_175 <= 0;
      findAndInsert_isFree_176 <= 0;
      findAndInsert_root_177 <= 0;
      findAndInsert_next_178 <= 0;
      findAndInsert_isLeaf_179 <= 0;
      findAndInsert_isFree_180 <= 0;
      findAndInsert_i_181 <= 0;
      findAndInsert_notFull_182 <= 0;
      findAndInsert_i_183 <= 0;
      findAndInsert_notFull_184 <= 0;
      findAndInsert_index_185 <= 0;
      findAndInsert_size_186 <= 0;
      findAndInsert_isLeaf_187 <= 0;
      findAndInsert_nextFree_188 <= 0;
      findAndInsert_Key_0_189 <= 0;
      findAndInsert_KeyCompares_0_190 <= 0;
      findAndInsert_KeyCollapse_0_191 <= 0;
      findAndInsert_Data_0_192 <= 0;
      findAndInsert_Key_1_193 <= 0;
      findAndInsert_KeyCompares_1_194 <= 0;
      findAndInsert_KeyCollapse_1_195 <= 0;
      findAndInsert_Data_1_196 <= 0;
      findAndInsert_Key_2_197 <= 0;
      findAndInsert_KeyCompares_2_198 <= 0;
      findAndInsert_KeyCollapse_2_199 <= 0;
      findAndInsert_Data_2_200 <= 0;
      findAndInsert_Key_3_201 <= 0;
      findAndInsert_KeyCompares_3_202 <= 0;
      findAndInsert_KeyCollapse_3_203 <= 0;
      findAndInsert_Data_3_204 <= 0;
      findAndInsert_Found_205 <= 0;
      findAndInsert_Key_206 <= 0;
      findAndInsert_FoundKey_207 <= 0;
      findAndInsert_Data_208 <= 0;
      findAndInsert_BtreeIndex_209 <= 0;
      findAndInsert_StuckIndex_210 <= 0;
      findAndInsert_MergeSuccess_211 <= 0;
      findAndInsert_index_212 <= 0;
      findAndInsert_size_213 <= 0;
      findAndInsert_isLeaf_214 <= 0;
      findAndInsert_nextFree_215 <= 0;
      findAndInsert_Key_0_216 <= 0;
      findAndInsert_KeyCompares_0_217 <= 0;
      findAndInsert_KeyCollapse_0_218 <= 0;
      findAndInsert_Data_0_219 <= 0;
      findAndInsert_Key_1_220 <= 0;
      findAndInsert_KeyCompares_1_221 <= 0;
      findAndInsert_KeyCollapse_1_222 <= 0;
      findAndInsert_Data_1_223 <= 0;
      findAndInsert_Key_2_224 <= 0;
      findAndInsert_KeyCompares_2_225 <= 0;
      findAndInsert_KeyCollapse_2_226 <= 0;
      findAndInsert_Data_2_227 <= 0;
      findAndInsert_Key_3_228 <= 0;
      findAndInsert_KeyCompares_3_229 <= 0;
      findAndInsert_KeyCollapse_3_230 <= 0;
      findAndInsert_Data_3_231 <= 0;
      findAndInsert_Found_232 <= 0;
      findAndInsert_Key_233 <= 0;
      findAndInsert_FoundKey_234 <= 0;
      findAndInsert_Data_235 <= 0;
      findAndInsert_BtreeIndex_236 <= 0;
      findAndInsert_StuckIndex_237 <= 0;
      findAndInsert_MergeSuccess_238 <= 0;
      findAndInsert_index_239 <= 0;
      findAndInsert_size_240 <= 0;
      findAndInsert_isLeaf_241 <= 0;
      findAndInsert_nextFree_242 <= 0;
      findAndInsert_Key_0_243 <= 0;
      findAndInsert_KeyCompares_0_244 <= 0;
      findAndInsert_KeyCollapse_0_245 <= 0;
      findAndInsert_Data_0_246 <= 0;
      findAndInsert_Key_1_247 <= 0;
      findAndInsert_KeyCompares_1_248 <= 0;
      findAndInsert_KeyCollapse_1_249 <= 0;
      findAndInsert_Data_1_250 <= 0;
      findAndInsert_Key_2_251 <= 0;
      findAndInsert_KeyCompares_2_252 <= 0;
      findAndInsert_KeyCollapse_2_253 <= 0;
      findAndInsert_Data_2_254 <= 0;
      findAndInsert_Key_3_255 <= 0;
      findAndInsert_KeyCompares_3_256 <= 0;
      findAndInsert_KeyCollapse_3_257 <= 0;
      findAndInsert_Data_3_258 <= 0;
      findAndInsert_Found_259 <= 0;
      findAndInsert_Key_260 <= 0;
      findAndInsert_FoundKey_261 <= 0;
      findAndInsert_Data_262 <= 0;
      findAndInsert_BtreeIndex_263 <= 0;
      findAndInsert_StuckIndex_264 <= 0;
      findAndInsert_MergeSuccess_265 <= 0;
      findAndInsert_childIndex_266 <= 0;
      findAndInsert_leftIndex_267 <= 0;
      findAndInsert_midKey_268 <= 0;
      findAndInsert_root_269 <= 0;
      findAndInsert_next_270 <= 0;
      findAndInsert_isLeaf_271 <= 0;
      findAndInsert_isFree_272 <= 0;
      findAndInsert_index_273 <= 0;
      findAndInsert_size_274 <= 0;
      findAndInsert_isLeaf_275 <= 0;
      findAndInsert_nextFree_276 <= 0;
      findAndInsert_Key_0_277 <= 0;
      findAndInsert_KeyCompares_0_278 <= 0;
      findAndInsert_KeyCollapse_0_279 <= 0;
      findAndInsert_Data_0_280 <= 0;
      findAndInsert_Key_1_281 <= 0;
      findAndInsert_KeyCompares_1_282 <= 0;
      findAndInsert_KeyCollapse_1_283 <= 0;
      findAndInsert_Data_1_284 <= 0;
      findAndInsert_Key_2_285 <= 0;
      findAndInsert_KeyCompares_2_286 <= 0;
      findAndInsert_KeyCollapse_2_287 <= 0;
      findAndInsert_Data_2_288 <= 0;
      findAndInsert_Key_3_289 <= 0;
      findAndInsert_KeyCompares_3_290 <= 0;
      findAndInsert_KeyCollapse_3_291 <= 0;
      findAndInsert_Data_3_292 <= 0;
      findAndInsert_Found_293 <= 0;
      findAndInsert_Key_294 <= 0;
      findAndInsert_FoundKey_295 <= 0;
      findAndInsert_Data_296 <= 0;
      findAndInsert_BtreeIndex_297 <= 0;
      findAndInsert_StuckIndex_298 <= 0;
      findAndInsert_MergeSuccess_299 <= 0;
      findAndInsert_index_300 <= 0;
      findAndInsert_size_301 <= 0;
      findAndInsert_isLeaf_302 <= 0;
      findAndInsert_nextFree_303 <= 0;
      findAndInsert_Key_0_304 <= 0;
      findAndInsert_KeyCompares_0_305 <= 0;
      findAndInsert_KeyCollapse_0_306 <= 0;
      findAndInsert_Data_0_307 <= 0;
      findAndInsert_Key_1_308 <= 0;
      findAndInsert_KeyCompares_1_309 <= 0;
      findAndInsert_KeyCollapse_1_310 <= 0;
      findAndInsert_Data_1_311 <= 0;
      findAndInsert_Key_2_312 <= 0;
      findAndInsert_KeyCompares_2_313 <= 0;
      findAndInsert_KeyCollapse_2_314 <= 0;
      findAndInsert_Data_2_315 <= 0;
      findAndInsert_Key_3_316 <= 0;
      findAndInsert_KeyCompares_3_317 <= 0;
      findAndInsert_KeyCollapse_3_318 <= 0;
      findAndInsert_Data_3_319 <= 0;
      findAndInsert_Found_320 <= 0;
      findAndInsert_Key_321 <= 0;
      findAndInsert_FoundKey_322 <= 0;
      findAndInsert_Data_323 <= 0;
      findAndInsert_BtreeIndex_324 <= 0;
      findAndInsert_StuckIndex_325 <= 0;
      findAndInsert_MergeSuccess_326 <= 0;
      findAndInsert_childKey_327 <= 0;
      findAndInsert_childData_328 <= 0;
      findAndInsert_indexLeft_329 <= 0;
      findAndInsert_indexRight_330 <= 0;
      findAndInsert_midKey_331 <= 0;
      findAndInsert_success_332 <= 0;
      findAndInsert_test_333 <= 0;
      findAndInsert_next_334 <= 0;
      findAndInsert_root_335 <= 0;
      findAndInsert_isFree_336 <= 0;
      stuckIsLeaf_7_requestedAt <= -1;
      stuckIsLeaf_8_requestedAt <= -1;
      stuckIsFree_11_requestedAt <= -1;
      freeNext_9_requestedAt <= -1;
      freeNext_10_requestedAt <= -1;
      stuckSize_5_requestedAt <= -1;
      stuckSize_6_requestedAt <= -1;
      stuckKeys_1_requestedAt <= -1;
      stuckKeys_2_requestedAt <= -1;
      stuckData_3_requestedAt <= -1;
      stuckData_4_requestedAt <= -1;
    end
    else if (processCurrent == 6) begin
      case(findAndInsert_pc)
        0: begin
          findAndInsert_k_45 <= 10;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        1: begin
          findAndInsert_d_46 <= 20;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        2: begin
          findAndInsert_BtreeIndex_73 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        3: begin
          findAndInsert_index_49 <= findAndInsert_BtreeIndex_73;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        4: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        5: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        6: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        7: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        8: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        9: begin
          findAndInsert_size_50 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_56 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_60 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_64 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_68 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        10: begin
          if (findAndInsert_isLeaf_51 == 0) begin
            findAndInsert_pc <= 17;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        11: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 == findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 == findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 == findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 == findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0803:<init>|  Btree.java:0802:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        12: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        13: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        14: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Key_70 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Key_70 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Key_70 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Key_70 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0846:<init>|  Btree.java:0845:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        15: begin
          findAndInsert_pc <= 23;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2260:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        16: begin
          findAndInsert_pc <= 23;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        17: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        18: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        19: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        20: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        21: begin
          findAndInsert_BtreeIndex_73 <= findAndInsert_Data_72;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:2264:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        22: begin
          findAndInsert_pc <= 3;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2265:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        23: begin
          if (findAndInsert_Found_69 == 0) begin
            findAndInsert_pc <= 26;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        24: begin
          if (findAndInsert_StuckIndex_74 == findAndInsert_size_50) begin
            findAndInsert_size_50 <= findAndInsert_size_50+1;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:2295:Then|  Chip.java:0606:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        25: begin
          findAndInsert_pc <= 37;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        26: begin
          findAndInsert_notFull_77 <= findAndInsert_size_50< 4 ? 1 : 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Lt|  Btree.java:2299:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        27: begin
          if (findAndInsert_notFull_77 == 0) begin
            findAndInsert_pc <= 36;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        28: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        29: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        30: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        31: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        32: begin
          findAndInsert_size_50 <= findAndInsert_size_50+1;
          if (3 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_3_65 <= findAndInsert_Key_2_61;
            findAndInsert_Data_3_68 <= findAndInsert_Data_2_64;
          end
          if (2 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_2_61 <= findAndInsert_Key_1_57;
            findAndInsert_Data_2_64 <= findAndInsert_Data_1_60;
          end
          if (1 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_1_57 <= findAndInsert_Key_0_53;
            findAndInsert_Data_1_60 <= findAndInsert_Data_0_56;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0702:<init>|  Btree.java:0701:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        33: begin
          findAndInsert_Found_69 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:2305:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        34: begin
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0588:<init>|  Chip.java:0587:COntinue|  Btree.java:2306:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        35: begin
          findAndInsert_pc <= 37;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        36: begin
          findAndInsert_pc <= 41;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2309:Else|  Chip.java:0616:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        37: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_49;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_50;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_49;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_53;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_57;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_61;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_65;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_49;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_56;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_60;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_64;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_68;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        38: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        39: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        40: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4172:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        41: begin
          findAndInsert_k_45 <= 20;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        42: begin
          findAndInsert_d_46 <= 30;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        43: begin
          findAndInsert_BtreeIndex_73 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        44: begin
          findAndInsert_index_49 <= findAndInsert_BtreeIndex_73;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        45: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        46: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        47: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        48: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        49: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        50: begin
          findAndInsert_size_50 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_56 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_60 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_64 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_68 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        51: begin
          if (findAndInsert_isLeaf_51 == 0) begin
            findAndInsert_pc <= 58;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        52: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 == findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 == findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 == findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 == findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0803:<init>|  Btree.java:0802:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        53: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        54: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        55: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Key_70 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Key_70 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Key_70 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Key_70 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0846:<init>|  Btree.java:0845:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        56: begin
          findAndInsert_pc <= 64;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2260:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        57: begin
          findAndInsert_pc <= 64;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        58: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        59: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        60: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        61: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        62: begin
          findAndInsert_BtreeIndex_73 <= findAndInsert_Data_72;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:2264:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        63: begin
          findAndInsert_pc <= 44;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2265:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        64: begin
          if (findAndInsert_Found_69 == 0) begin
            findAndInsert_pc <= 67;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        65: begin
          if (findAndInsert_StuckIndex_74 == findAndInsert_size_50) begin
            findAndInsert_size_50 <= findAndInsert_size_50+1;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:2295:Then|  Chip.java:0606:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        66: begin
          findAndInsert_pc <= 78;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        67: begin
          findAndInsert_notFull_79 <= findAndInsert_size_50< 4 ? 1 : 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Lt|  Btree.java:2299:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        68: begin
          if (findAndInsert_notFull_79 == 0) begin
            findAndInsert_pc <= 77;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        69: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        70: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        71: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        72: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        73: begin
          findAndInsert_size_50 <= findAndInsert_size_50+1;
          if (3 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_3_65 <= findAndInsert_Key_2_61;
            findAndInsert_Data_3_68 <= findAndInsert_Data_2_64;
          end
          if (2 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_2_61 <= findAndInsert_Key_1_57;
            findAndInsert_Data_2_64 <= findAndInsert_Data_1_60;
          end
          if (1 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_1_57 <= findAndInsert_Key_0_53;
            findAndInsert_Data_1_60 <= findAndInsert_Data_0_56;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0702:<init>|  Btree.java:0701:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        74: begin
          findAndInsert_Found_69 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:2305:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        75: begin
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0588:<init>|  Chip.java:0587:COntinue|  Btree.java:2306:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        76: begin
          findAndInsert_pc <= 78;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        77: begin
          findAndInsert_pc <= 82;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2309:Else|  Chip.java:0616:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        78: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_49;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_50;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_49;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_53;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_57;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_61;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_65;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_49;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_56;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_60;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_64;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_68;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        79: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        80: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        81: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4173:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        82: begin
          findAndInsert_k_45 <= 40;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        83: begin
          findAndInsert_d_46 <= 50;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        84: begin
          findAndInsert_BtreeIndex_73 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        85: begin
          findAndInsert_index_49 <= findAndInsert_BtreeIndex_73;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        86: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        87: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        88: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        89: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        90: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        91: begin
          findAndInsert_size_50 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_56 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_60 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_64 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_68 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        92: begin
          if (findAndInsert_isLeaf_51 == 0) begin
            findAndInsert_pc <= 99;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        93: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 == findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 == findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 == findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 == findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0803:<init>|  Btree.java:0802:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        94: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        95: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        96: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Key_70 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Key_70 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Key_70 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Key_70 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0846:<init>|  Btree.java:0845:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        97: begin
          findAndInsert_pc <= 105;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2260:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        98: begin
          findAndInsert_pc <= 105;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        99: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        100: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        101: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        102: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        103: begin
          findAndInsert_BtreeIndex_73 <= findAndInsert_Data_72;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:2264:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        104: begin
          findAndInsert_pc <= 85;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2265:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        105: begin
          if (findAndInsert_Found_69 == 0) begin
            findAndInsert_pc <= 108;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        106: begin
          if (findAndInsert_StuckIndex_74 == findAndInsert_size_50) begin
            findAndInsert_size_50 <= findAndInsert_size_50+1;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:2295:Then|  Chip.java:0606:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        107: begin
          findAndInsert_pc <= 119;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        108: begin
          findAndInsert_notFull_81 <= findAndInsert_size_50< 4 ? 1 : 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Lt|  Btree.java:2299:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        109: begin
          if (findAndInsert_notFull_81 == 0) begin
            findAndInsert_pc <= 118;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        110: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        111: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        112: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        113: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        114: begin
          findAndInsert_size_50 <= findAndInsert_size_50+1;
          if (3 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_3_65 <= findAndInsert_Key_2_61;
            findAndInsert_Data_3_68 <= findAndInsert_Data_2_64;
          end
          if (2 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_2_61 <= findAndInsert_Key_1_57;
            findAndInsert_Data_2_64 <= findAndInsert_Data_1_60;
          end
          if (1 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_1_57 <= findAndInsert_Key_0_53;
            findAndInsert_Data_1_60 <= findAndInsert_Data_0_56;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0702:<init>|  Btree.java:0701:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        115: begin
          findAndInsert_Found_69 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:2305:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        116: begin
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0588:<init>|  Chip.java:0587:COntinue|  Btree.java:2306:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        117: begin
          findAndInsert_pc <= 119;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        118: begin
          findAndInsert_pc <= 123;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2309:Else|  Chip.java:0616:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        119: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_49;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_50;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_49;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_53;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_57;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_61;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_65;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_49;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_56;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_60;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_64;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_68;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        120: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        121: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        122: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4174:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        123: begin
          findAndInsert_k_45 <= 30;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        124: begin
          findAndInsert_d_46 <= 40;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        125: begin
          findAndInsert_BtreeIndex_73 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        126: begin
          findAndInsert_index_49 <= findAndInsert_BtreeIndex_73;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        127: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        128: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        129: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        130: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        131: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        132: begin
          findAndInsert_size_50 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_56 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_60 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_64 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_68 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        133: begin
          if (findAndInsert_isLeaf_51 == 0) begin
            findAndInsert_pc <= 140;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        134: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 == findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 == findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 == findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 == findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0803:<init>|  Btree.java:0802:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        135: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        136: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        137: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Key_70 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Key_70 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Key_70 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Key_70 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0846:<init>|  Btree.java:0845:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        138: begin
          findAndInsert_pc <= 146;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2260:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        139: begin
          findAndInsert_pc <= 146;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        140: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        141: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        142: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        143: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        144: begin
          findAndInsert_BtreeIndex_73 <= findAndInsert_Data_72;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:2264:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        145: begin
          findAndInsert_pc <= 126;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2265:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        146: begin
          if (findAndInsert_Found_69 == 0) begin
            findAndInsert_pc <= 149;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        147: begin
          if (findAndInsert_StuckIndex_74 == findAndInsert_size_50) begin
            findAndInsert_size_50 <= findAndInsert_size_50+1;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:2295:Then|  Chip.java:0606:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        148: begin
          findAndInsert_pc <= 160;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        149: begin
          findAndInsert_notFull_83 <= findAndInsert_size_50< 4 ? 1 : 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Lt|  Btree.java:2299:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        150: begin
          if (findAndInsert_notFull_83 == 0) begin
            findAndInsert_pc <= 159;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        151: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        152: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        153: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        154: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        155: begin
          findAndInsert_size_50 <= findAndInsert_size_50+1;
          if (3 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_3_65 <= findAndInsert_Key_2_61;
            findAndInsert_Data_3_68 <= findAndInsert_Data_2_64;
          end
          if (2 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_2_61 <= findAndInsert_Key_1_57;
            findAndInsert_Data_2_64 <= findAndInsert_Data_1_60;
          end
          if (1 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_1_57 <= findAndInsert_Key_0_53;
            findAndInsert_Data_1_60 <= findAndInsert_Data_0_56;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0702:<init>|  Btree.java:0701:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        156: begin
          findAndInsert_Found_69 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:2305:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        157: begin
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0588:<init>|  Chip.java:0587:COntinue|  Btree.java:2306:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        158: begin
          findAndInsert_pc <= 160;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        159: begin
          findAndInsert_pc <= 164;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2309:Else|  Chip.java:0616:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        160: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_49;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_50;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_49;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_53;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_57;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_61;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_65;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_49;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_56;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_60;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_64;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_68;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        161: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        162: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        163: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4175:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        164: begin
          findAndInsert_index_84 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        165: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_84;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_84;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_84;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_84;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0269:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        166: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0269:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        167: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0269:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        168: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0269:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        169: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0269:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        170: begin
          findAndInsert_size_85 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_86 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_88 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_91 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_92 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_95 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_96 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_99 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_100 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_103 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0269:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        171: begin
          if (findAndInsert_size_85 < 4) begin
            findAndInsert_pc <= 217;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1532:<init>|  Btree.java:1531:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        172: begin
          findAndInsert_Key_0_115 <= findAndInsert_Key_0_88;
          findAndInsert_Data_0_118 <= findAndInsert_Data_0_91;
          findAndInsert_Key_1_119 <= findAndInsert_Key_1_92;
          findAndInsert_Data_1_122 <= findAndInsert_Data_1_95;
          findAndInsert_size_112 <= 2;
          findAndInsert_Key_0_142 <= findAndInsert_Key_2_96;
          findAndInsert_Data_0_145 <= findAndInsert_Data_2_99;
          findAndInsert_Key_1_146 <= findAndInsert_Key_3_100;
          findAndInsert_Data_1_149 <= findAndInsert_Data_3_103;
          findAndInsert_size_139 <= 2;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:1043:<init>|  Btree.java:1042:splitIntoTwo|  Btree.java:1549:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        173: begin
          findAndInsert_root_173 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:0077:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        174: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_root_173;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1278:<init>|  Chip.java:1277:ExecuteTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        175: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0079:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        176: begin
          findAndInsert_indexLeft_165 <= freeNext_freeNext_9_result_0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0080:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        177: begin
          if (findAndInsert_indexLeft_165 == 0) begin
            findAndInsert_returnCode <= 20;
            findAndInsert_stop <= 1;
          end
          findAndInsert_isLeaf_175 <= 1;
          findAndInsert_isFree_176 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0083:<init>|  Btree.java:0082:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        178: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_indexLeft_165;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_8_index_36 <= findAndInsert_indexLeft_165;
          findAndInsert_stuckIsLeaf_8_value_37 <= findAndInsert_isLeaf_175;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          findAndInsert_stuckIsFree_11_index_171 <= findAndInsert_indexLeft_165;
          findAndInsert_stuckIsFree_11_value_172 <= findAndInsert_isFree_176;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0098:<init>|  Btree.java:0097:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        179: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0110:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        180: begin
          findAndInsert_next_174 <= freeNext_freeNext_9_result_0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0111:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        181: begin
          findAndInsert_freeNext_10_index_169 <= findAndInsert_root_173;
          findAndInsert_freeNext_10_value_170 <= findAndInsert_next_174;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1341:<init>|  Chip.java:1340:ExecuteTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        182: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        183: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        184: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0115:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        185: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_indexLeft_165;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_112;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_indexLeft_165;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_115;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_119;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_123;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_127;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_indexLeft_165;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_118;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_122;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_126;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_130;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        186: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        187: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        188: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1551:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        189: begin
          findAndInsert_root_177 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:0077:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        190: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_root_177;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1278:<init>|  Chip.java:1277:ExecuteTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        191: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0079:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        192: begin
          findAndInsert_indexRight_166 <= freeNext_freeNext_9_result_0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0080:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        193: begin
          if (findAndInsert_indexRight_166 == 0) begin
            findAndInsert_returnCode <= 20;
            findAndInsert_stop <= 1;
          end
          findAndInsert_isLeaf_179 <= 1;
          findAndInsert_isFree_180 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0083:<init>|  Btree.java:0082:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        194: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_indexRight_166;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_8_index_36 <= findAndInsert_indexRight_166;
          findAndInsert_stuckIsLeaf_8_value_37 <= findAndInsert_isLeaf_179;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          findAndInsert_stuckIsFree_11_index_171 <= findAndInsert_indexRight_166;
          findAndInsert_stuckIsFree_11_value_172 <= findAndInsert_isFree_180;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0098:<init>|  Btree.java:0097:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        195: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0110:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        196: begin
          findAndInsert_next_178 <= freeNext_freeNext_9_result_0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0111:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        197: begin
          findAndInsert_freeNext_10_index_169 <= findAndInsert_root_177;
          findAndInsert_freeNext_10_value_170 <= findAndInsert_next_178;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1341:<init>|  Chip.java:1340:ExecuteTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        198: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        199: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        200: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0115:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        201: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_indexRight_166;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_139;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_indexRight_166;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_142;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_146;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_150;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_154;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_indexRight_166;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_145;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_149;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_153;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_157;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        202: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        203: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        204: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1552:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        205: begin
          case (findAndInsert_size_112)
            1: begin
              findAndInsert_Key_132 <= findAndInsert_Key_0_115;
              findAndInsert_Data_134 <= findAndInsert_Data_0_118;
            end
            2: begin
              findAndInsert_Key_132 <= findAndInsert_Key_1_119;
              findAndInsert_Data_134 <= findAndInsert_Data_1_122;
            end
            3: begin
              findAndInsert_Key_132 <= findAndInsert_Key_2_123;
              findAndInsert_Data_134 <= findAndInsert_Data_2_126;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0532:<init>|  Btree.java:0531:LastElement|  Btree.java:1554:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        206: begin
          findAndInsert_Key_159 <= findAndInsert_Key_0_142;
          findAndInsert_Data_161 <= findAndInsert_Data_0_145;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0505:<init>|  Btree.java:0504:FirstElement|  Btree.java:1555:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        207: begin
          findAndInsert_midKey_167 <= (findAndInsert_Key_132 + findAndInsert_Key_159) / 2;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0829:<init>|  Chip.java:0828:Average|  Btree.java:1556:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        208: begin
          findAndInsert_size_85 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0396:<init>|  Btree.java:0395:Clear|  Btree.java:1557:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        209: begin
          case (findAndInsert_size_85)
            0: begin
              findAndInsert_Key_0_88 <= findAndInsert_midKey_167;
              findAndInsert_Data_0_91 <= findAndInsert_indexLeft_165;
            end
            1: begin
              findAndInsert_Key_1_92 <= findAndInsert_midKey_167;
              findAndInsert_Data_1_95 <= findAndInsert_indexLeft_165;
            end
            2: begin
              findAndInsert_Key_2_96 <= findAndInsert_midKey_167;
              findAndInsert_Data_2_99 <= findAndInsert_indexLeft_165;
            end
            3: begin
              findAndInsert_Key_3_100 <= findAndInsert_midKey_167;
              findAndInsert_Data_3_103 <= findAndInsert_indexLeft_165;
            end
          endcase
          findAndInsert_size_85 <= findAndInsert_size_85+1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0425:<init>|  Btree.java:0424:Push|  Btree.java:1558:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        210: begin
          case (findAndInsert_size_85)
            0: begin
              findAndInsert_Key_0_88 <= findAndInsert_midKey_167;
              findAndInsert_Data_0_91 <= findAndInsert_indexRight_166;
            end
            1: begin
              findAndInsert_Key_1_92 <= findAndInsert_midKey_167;
              findAndInsert_Data_1_95 <= findAndInsert_indexRight_166;
            end
            2: begin
              findAndInsert_Key_2_96 <= findAndInsert_midKey_167;
              findAndInsert_Data_2_99 <= findAndInsert_indexRight_166;
            end
            3: begin
              findAndInsert_Key_3_100 <= findAndInsert_midKey_167;
              findAndInsert_Data_3_103 <= findAndInsert_indexRight_166;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0482:<init>|  Btree.java:0481:SetPastLastElement|  Btree.java:1559:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        211: begin
          findAndInsert_isLeaf_86 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:1560:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        212: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_84;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_85;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_8_index_36 <= findAndInsert_index_84;
          findAndInsert_stuckIsLeaf_8_value_37 <= findAndInsert_isLeaf_86;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_84;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_88;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_92;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_96;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_100;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_84;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_91;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_95;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_99;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_103;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:1561:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        213: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:1561:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        214: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:1561:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        215: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:1561:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        216: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:1561:code|  Chip.java:0526:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:4177:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        217: begin
          findAndInsert_k_45 <= 50;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        218: begin
          findAndInsert_d_46 <= 60;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        219: begin
          findAndInsert_BtreeIndex_73 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        220: begin
          findAndInsert_index_49 <= findAndInsert_BtreeIndex_73;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        221: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        222: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        223: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        224: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        225: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        226: begin
          findAndInsert_size_50 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_56 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_60 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_64 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_68 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        227: begin
          if (findAndInsert_isLeaf_51 == 0) begin
            findAndInsert_pc <= 234;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        228: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 == findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 == findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 == findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 == findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0803:<init>|  Btree.java:0802:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        229: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        230: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        231: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Key_70 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Key_70 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Key_70 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Key_70 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0846:<init>|  Btree.java:0845:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        232: begin
          findAndInsert_pc <= 240;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2260:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        233: begin
          findAndInsert_pc <= 240;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        234: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        235: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        236: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        237: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        238: begin
          findAndInsert_BtreeIndex_73 <= findAndInsert_Data_72;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:2264:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        239: begin
          findAndInsert_pc <= 220;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2265:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        240: begin
          if (findAndInsert_Found_69 == 0) begin
            findAndInsert_pc <= 243;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        241: begin
          if (findAndInsert_StuckIndex_74 == findAndInsert_size_50) begin
            findAndInsert_size_50 <= findAndInsert_size_50+1;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:2295:Then|  Chip.java:0606:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        242: begin
          findAndInsert_pc <= 254;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        243: begin
          findAndInsert_notFull_182 <= findAndInsert_size_50< 4 ? 1 : 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Lt|  Btree.java:2299:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        244: begin
          if (findAndInsert_notFull_182 == 0) begin
            findAndInsert_pc <= 253;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        245: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        246: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        247: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        248: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        249: begin
          findAndInsert_size_50 <= findAndInsert_size_50+1;
          if (3 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_3_65 <= findAndInsert_Key_2_61;
            findAndInsert_Data_3_68 <= findAndInsert_Data_2_64;
          end
          if (2 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_2_61 <= findAndInsert_Key_1_57;
            findAndInsert_Data_2_64 <= findAndInsert_Data_1_60;
          end
          if (1 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_1_57 <= findAndInsert_Key_0_53;
            findAndInsert_Data_1_60 <= findAndInsert_Data_0_56;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0702:<init>|  Btree.java:0701:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        250: begin
          findAndInsert_Found_69 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:2305:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        251: begin
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0588:<init>|  Chip.java:0587:COntinue|  Btree.java:2306:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        252: begin
          findAndInsert_pc <= 254;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        253: begin
          findAndInsert_pc <= 258;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2309:Else|  Chip.java:0616:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        254: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_49;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_50;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_49;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_53;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_57;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_61;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_65;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_49;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_56;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_60;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_64;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_68;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        255: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        256: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        257: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4179:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        258: begin
          findAndInsert_k_45 <= 60;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        259: begin
          findAndInsert_d_46 <= 70;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        260: begin
          findAndInsert_BtreeIndex_73 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        261: begin
          findAndInsert_index_49 <= findAndInsert_BtreeIndex_73;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        262: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        263: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        264: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        265: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        266: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        267: begin
          findAndInsert_size_50 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_56 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_60 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_64 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_68 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:2256:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        268: begin
          if (findAndInsert_isLeaf_51 == 0) begin
            findAndInsert_pc <= 275;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        269: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 == findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 == findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 == findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 == findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0803:<init>|  Btree.java:0802:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        270: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        271: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0824:<init>|  Btree.java:0823:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        272: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Key_70 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Key_70 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Key_70 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Key_70 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0846:<init>|  Btree.java:0845:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        273: begin
          findAndInsert_pc <= 281;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2260:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        274: begin
          findAndInsert_pc <= 281;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        275: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        276: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        277: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        278: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        279: begin
          findAndInsert_BtreeIndex_73 <= findAndInsert_Data_72;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:2264:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        280: begin
          findAndInsert_pc <= 261;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2265:Branch|  Btree.java:1415:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0526:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        281: begin
          if (findAndInsert_Found_69 == 0) begin
            findAndInsert_pc <= 284;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        282: begin
          if (findAndInsert_StuckIndex_74 == findAndInsert_size_50) begin
            findAndInsert_size_50 <= findAndInsert_size_50+1;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:2295:Then|  Chip.java:0606:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        283: begin
          findAndInsert_pc <= 295;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        284: begin
          findAndInsert_notFull_184 <= findAndInsert_size_50< 4 ? 1 : 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Lt|  Btree.java:2299:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        285: begin
          if (findAndInsert_notFull_184 == 0) begin
            findAndInsert_pc <= 294;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        286: begin
          findAndInsert_KeyCompares_0_54 <= findAndInsert_k_45 <= findAndInsert_Key_0_53 && 0 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_0_55 <= 0;
          findAndInsert_KeyCompares_1_58 <= findAndInsert_k_45 >  findAndInsert_Key_0_53 && findAndInsert_k_45 <= findAndInsert_Key_1_57 && 1 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_1_59 <= 1;
          findAndInsert_KeyCompares_2_62 <= findAndInsert_k_45 >  findAndInsert_Key_1_57 && findAndInsert_k_45 <= findAndInsert_Key_2_61 && 2 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_2_63 <= 2;
          findAndInsert_KeyCompares_3_66 <= findAndInsert_k_45 >  findAndInsert_Key_2_61 && findAndInsert_k_45 <= findAndInsert_Key_3_65 && 3 < findAndInsert_size_50;
          findAndInsert_KeyCollapse_3_67 <= 3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0939:<init>|  Btree.java:0938:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        287: begin
          if (findAndInsert_KeyCompares_1_58) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_1_59;
          end
          if (findAndInsert_KeyCompares_3_66) begin
            findAndInsert_KeyCompares_2_62 <= 1;
            findAndInsert_KeyCollapse_2_63 <= findAndInsert_KeyCollapse_3_67;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        288: begin
          if (findAndInsert_KeyCompares_2_62) begin
            findAndInsert_KeyCompares_0_54 <= 1;
            findAndInsert_KeyCollapse_0_55 <= findAndInsert_KeyCollapse_2_63;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0975:<init>|  Btree.java:0974:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        289: begin
          if (findAndInsert_KeyCompares_0_54) begin
            findAndInsert_Found_69 <= 1;
            case (findAndInsert_KeyCollapse_0_55)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_0_53;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_1_57;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_2_61;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_FoundKey_71 <= findAndInsert_Key_3_65;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          else begin
            findAndInsert_Found_69 <= 0;
            case (findAndInsert_size_50)
              0: begin
                findAndInsert_StuckIndex_74 <= 0;
                findAndInsert_Data_72 <= findAndInsert_Data_0_56;
              end
              1: begin
                findAndInsert_StuckIndex_74 <= 1;
                findAndInsert_Data_72 <= findAndInsert_Data_1_60;
              end
              2: begin
                findAndInsert_StuckIndex_74 <= 2;
                findAndInsert_Data_72 <= findAndInsert_Data_2_64;
              end
              3: begin
                findAndInsert_StuckIndex_74 <= 3;
                findAndInsert_Data_72 <= findAndInsert_Data_3_68;
              end
            endcase
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0997:<init>|  Btree.java:0996:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        290: begin
          findAndInsert_size_50 <= findAndInsert_size_50+1;
          if (3 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_3_65 <= findAndInsert_Key_2_61;
            findAndInsert_Data_3_68 <= findAndInsert_Data_2_64;
          end
          if (2 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_2_61 <= findAndInsert_Key_1_57;
            findAndInsert_Data_2_64 <= findAndInsert_Data_1_60;
          end
          if (1 > findAndInsert_StuckIndex_74) begin
            findAndInsert_Key_1_57 <= findAndInsert_Key_0_53;
            findAndInsert_Data_1_60 <= findAndInsert_Data_0_56;
          end
          case (findAndInsert_StuckIndex_74)
            0: begin
              findAndInsert_Key_0_53 <= findAndInsert_k_45;
              findAndInsert_Data_0_56 <= findAndInsert_d_46;
            end
            1: begin
              findAndInsert_Key_1_57 <= findAndInsert_k_45;
              findAndInsert_Data_1_60 <= findAndInsert_d_46;
            end
            2: begin
              findAndInsert_Key_2_61 <= findAndInsert_k_45;
              findAndInsert_Data_2_64 <= findAndInsert_d_46;
            end
            3: begin
              findAndInsert_Key_3_65 <= findAndInsert_k_45;
              findAndInsert_Data_3_68 <= findAndInsert_d_46;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0702:<init>|  Btree.java:0701:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        291: begin
          findAndInsert_Found_69 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:2305:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        292: begin
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0588:<init>|  Chip.java:0587:COntinue|  Btree.java:2306:Then|  Chip.java:0606:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        293: begin
          findAndInsert_pc <= 295;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        294: begin
          findAndInsert_pc <= 299;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:2309:Else|  Chip.java:0616:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0616:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        295: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_49;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_50;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_49;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_53;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_57;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_61;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_65;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_49;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_56;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_60;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_64;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_68;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        296: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        297: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        298: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0338:stuckPut|  Btree.java:2314:code|  Chip.java:0526:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:4180:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        299: begin
          findAndInsert_i_47 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4182:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        300: begin
          findAndInsert_index_185 <= findAndInsert_i_47;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        301: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_185;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_185;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_185;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_185;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        302: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        303: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        304: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        305: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        306: begin
          findAndInsert_size_186 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_187 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_189 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_192 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_193 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_196 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_197 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_200 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_201 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_204 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        307: begin
          case (findAndInsert_size_186)
            0: begin
              findAndInsert_Key_206 <= findAndInsert_Key_0_189;
              findAndInsert_Data_208 <= findAndInsert_Data_0_192;
            end
            1: begin
              findAndInsert_Key_206 <= findAndInsert_Key_1_193;
              findAndInsert_Data_208 <= findAndInsert_Data_1_196;
            end
            2: begin
              findAndInsert_Key_206 <= findAndInsert_Key_2_197;
              findAndInsert_Data_208 <= findAndInsert_Data_2_200;
            end
            3: begin
              findAndInsert_Key_206 <= findAndInsert_Key_3_201;
              findAndInsert_Data_208 <= findAndInsert_Data_3_204;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0559:<init>|  Btree.java:0558:PastLastElement|  Btree.java:1655:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        308: begin
          findAndInsert_childIndex_266 <= findAndInsert_Data_208;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:1656:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        309: begin
          findAndInsert_index_212 <= findAndInsert_childIndex_266;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        310: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_212;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_212;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_212;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_212;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        311: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        312: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        313: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        314: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        315: begin
          findAndInsert_size_213 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_214 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_216 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_219 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_220 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_223 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_224 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_227 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_228 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_231 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        316: begin
          
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:1660:<init>|  Btree.java:1659:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        317: begin
          findAndInsert_Key_0_243 <= findAndInsert_Key_0_216;
          findAndInsert_Data_0_246 <= findAndInsert_Data_0_219;
          findAndInsert_Key_1_247 <= findAndInsert_Key_1_220;
          findAndInsert_Data_1_250 <= findAndInsert_Data_1_223;
          findAndInsert_size_240 <= 2;
          findAndInsert_Key_0_216 <= findAndInsert_Key_2_224;
          findAndInsert_Data_0_219 <= findAndInsert_Data_2_227;
          findAndInsert_Key_1_220 <= findAndInsert_Key_3_228;
          findAndInsert_Data_1_223 <= findAndInsert_Data_3_231;
          findAndInsert_size_213 <= 2;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:1126:<init>|  Btree.java:1125:splitLow|  Btree.java:1669:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        318: begin
          findAndInsert_root_269 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:0077:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        319: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_root_269;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1278:<init>|  Chip.java:1277:ExecuteTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        320: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0079:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        321: begin
          findAndInsert_leftIndex_267 <= freeNext_freeNext_9_result_0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0080:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        322: begin
          if (findAndInsert_leftIndex_267 == 0) begin
            findAndInsert_returnCode <= 20;
            findAndInsert_stop <= 1;
          end
          findAndInsert_isLeaf_271 <= 1;
          findAndInsert_isFree_272 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0083:<init>|  Btree.java:0082:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        323: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_leftIndex_267;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_8_index_36 <= findAndInsert_leftIndex_267;
          findAndInsert_stuckIsLeaf_8_value_37 <= findAndInsert_isLeaf_271;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          findAndInsert_stuckIsFree_11_index_171 <= findAndInsert_leftIndex_267;
          findAndInsert_stuckIsFree_11_value_172 <= findAndInsert_isFree_272;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0098:<init>|  Btree.java:0097:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        324: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0110:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        325: begin
          findAndInsert_next_270 <= freeNext_freeNext_9_result_0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0111:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        326: begin
          findAndInsert_freeNext_10_index_169 <= findAndInsert_root_269;
          findAndInsert_freeNext_10_value_170 <= findAndInsert_next_270;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1341:<init>|  Chip.java:1340:ExecuteTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        327: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        328: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        329: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0115:allocate|  Btree.java:0152:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        330: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_leftIndex_267;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_240;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_leftIndex_267;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_243;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_247;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_251;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_255;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_leftIndex_267;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_246;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_250;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_254;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_258;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        331: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        332: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        333: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        334: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_childIndex_266;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_213;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_childIndex_266;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_216;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_220;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_224;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_228;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_childIndex_266;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_219;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_223;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_227;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_231;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        335: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        336: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        337: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        338: begin
          case (findAndInsert_size_240)
            1: begin
              findAndInsert_Key_260 <= findAndInsert_Key_0_243;
              findAndInsert_Data_262 <= findAndInsert_Data_0_246;
            end
            2: begin
              findAndInsert_Key_260 <= findAndInsert_Key_1_247;
              findAndInsert_Data_262 <= findAndInsert_Data_1_250;
            end
            3: begin
              findAndInsert_Key_260 <= findAndInsert_Key_2_251;
              findAndInsert_Data_262 <= findAndInsert_Data_2_254;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0532:<init>|  Btree.java:0531:LastElement|  Btree.java:1672:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        339: begin
          findAndInsert_Key_233 <= findAndInsert_Key_0_216;
          findAndInsert_Data_235 <= findAndInsert_Data_0_219;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0505:<init>|  Btree.java:0504:FirstElement|  Btree.java:1673:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        340: begin
          findAndInsert_midKey_268 <= (findAndInsert_Key_260 + findAndInsert_Key_233) / 2;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0829:<init>|  Chip.java:0828:Average|  Btree.java:1674:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        341: begin
          case (findAndInsert_size_186)
            0: begin
              findAndInsert_Key_0_189 <= findAndInsert_midKey_268;
              findAndInsert_Data_0_192 <= findAndInsert_leftIndex_267;
            end
            1: begin
              findAndInsert_Key_1_193 <= findAndInsert_midKey_268;
              findAndInsert_Data_1_196 <= findAndInsert_leftIndex_267;
            end
            2: begin
              findAndInsert_Key_2_197 <= findAndInsert_midKey_268;
              findAndInsert_Data_2_200 <= findAndInsert_leftIndex_267;
            end
            3: begin
              findAndInsert_Key_3_201 <= findAndInsert_midKey_268;
              findAndInsert_Data_3_204 <= findAndInsert_leftIndex_267;
            end
          endcase
          findAndInsert_size_186 <= findAndInsert_size_186+1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0425:<init>|  Btree.java:0424:Push|  Btree.java:1675:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        342: begin
          case (findAndInsert_size_186)
            0: begin
              findAndInsert_Key_0_189 <= findAndInsert_midKey_268;
              findAndInsert_Data_0_192 <= findAndInsert_childIndex_266;
            end
            1: begin
              findAndInsert_Key_1_193 <= findAndInsert_midKey_268;
              findAndInsert_Data_1_196 <= findAndInsert_childIndex_266;
            end
            2: begin
              findAndInsert_Key_2_197 <= findAndInsert_midKey_268;
              findAndInsert_Data_2_200 <= findAndInsert_childIndex_266;
            end
            3: begin
              findAndInsert_Key_3_201 <= findAndInsert_midKey_268;
              findAndInsert_Data_3_204 <= findAndInsert_childIndex_266;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0482:<init>|  Btree.java:0481:SetPastLastElement|  Btree.java:1676:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        343: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_185;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_186;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_185;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_189;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_193;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_197;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_201;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_185;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_192;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_196;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_200;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_204;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        344: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        345: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        346: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:4183:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        347: begin
          findAndInsert_i_47 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4185:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        348: begin
          findAndInsert_j_48 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0672:<init>|  Chip.java:0671:RegisterSet|  Btree.java:4185:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        349: begin
          findAndInsert_index_0 <= findAndInsert_i_47;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        350: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_0;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_0;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_0;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_0;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        351: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        352: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        353: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        354: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        355: begin
          findAndInsert_size_1 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_2 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_4 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_7 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_8 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_11 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_12 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_15 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_16 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_19 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:4186:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        356: begin
          if (findAndInsert_i_47 == 0 && findAndInsert_size_1 > 1) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          else begin
            if (findAndInsert_i_47 == 0 || findAndInsert_size_1 < 1) begin
              findAndInsert_pc <= 400;
            end
            else begin
              findAndInsert_pc <= findAndInsert_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1770:<init>|  Btree.java:1769:mergePermitted|  Btree.java:1878:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        357: begin
          case (findAndInsert_j_48)
            0: begin
              findAndInsert_indexLeft_329 <= findAndInsert_Data_0_7;
              findAndInsert_indexRight_330 <= findAndInsert_Data_1_11;
            end
            1: begin
              findAndInsert_indexLeft_329 <= findAndInsert_Data_1_11;
              findAndInsert_indexRight_330 <= findAndInsert_Data_2_15;
            end
            2: begin
              findAndInsert_indexLeft_329 <= findAndInsert_Data_2_15;
              findAndInsert_indexRight_330 <= findAndInsert_Data_3_19;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:1881:<init>|  Btree.java:1880:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        358: begin
          findAndInsert_index_273 <= findAndInsert_indexLeft_329;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        359: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_273;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_273;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_273;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_273;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        360: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        361: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        362: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        363: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        364: begin
          findAndInsert_size_274 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_275 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_277 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_280 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_281 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_284 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_285 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_288 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_289 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_292 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1895:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        365: begin
          findAndInsert_index_300 <= findAndInsert_indexRight_330;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0693:<init>|  Chip.java:0692:Copy|  Btree.java:0263:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        366: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_300;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_300;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_300;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_300;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0274:<init>|  Btree.java:0273:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        367: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        368: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        369: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        370: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0291:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        371: begin
          findAndInsert_size_301 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_302 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_304 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_307 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_308 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_311 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_312 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_315 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_316 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_319 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0294:<init>|  Btree.java:0293:stuckGet|  Btree.java:0264:stuckGet|  Btree.java:1896:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        372: begin
          if (findAndInsert_isLeaf_275 == 0) begin
            findAndInsert_pc <= 400;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        373: begin
          if (findAndInsert_isLeaf_302 == 0) begin
            findAndInsert_pc <= 399;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1396:<init>|  Btree.java:1395:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        374: begin
          findAndInsert_MergeSuccess_299 <= 0;
          case (findAndInsert_size_274)
            0: begin
              case (findAndInsert_size_301)
                0: begin
                  findAndInsert_size_274 <= findAndInsert_size_274 + 0;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                1: begin
                  findAndInsert_Key_0_277 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_0_280 <= findAndInsert_Data_0_307;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 1;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                2: begin
                  findAndInsert_Key_0_277 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_0_280 <= findAndInsert_Data_0_307;
                  findAndInsert_Key_1_281 <= findAndInsert_Key_1_308;
                  findAndInsert_Data_1_284 <= findAndInsert_Data_1_311;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 2;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                3: begin
                  findAndInsert_Key_0_277 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_0_280 <= findAndInsert_Data_0_307;
                  findAndInsert_Key_1_281 <= findAndInsert_Key_1_308;
                  findAndInsert_Data_1_284 <= findAndInsert_Data_1_311;
                  findAndInsert_Key_2_285 <= findAndInsert_Key_2_312;
                  findAndInsert_Data_2_288 <= findAndInsert_Data_2_315;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 3;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                4: begin
                  findAndInsert_Key_0_277 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_0_280 <= findAndInsert_Data_0_307;
                  findAndInsert_Key_1_281 <= findAndInsert_Key_1_308;
                  findAndInsert_Data_1_284 <= findAndInsert_Data_1_311;
                  findAndInsert_Key_2_285 <= findAndInsert_Key_2_312;
                  findAndInsert_Data_2_288 <= findAndInsert_Data_2_315;
                  findAndInsert_Key_3_289 <= findAndInsert_Key_3_316;
                  findAndInsert_Data_3_292 <= findAndInsert_Data_3_319;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 4;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
              endcase
            end
            1: begin
              case (findAndInsert_size_301)
                0: begin
                  findAndInsert_size_274 <= findAndInsert_size_274 + 0;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                1: begin
                  findAndInsert_Key_1_281 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_1_284 <= findAndInsert_Data_0_307;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 1;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                2: begin
                  findAndInsert_Key_1_281 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_1_284 <= findAndInsert_Data_0_307;
                  findAndInsert_Key_2_285 <= findAndInsert_Key_1_308;
                  findAndInsert_Data_2_288 <= findAndInsert_Data_1_311;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 2;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                3: begin
                  findAndInsert_Key_1_281 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_1_284 <= findAndInsert_Data_0_307;
                  findAndInsert_Key_2_285 <= findAndInsert_Key_1_308;
                  findAndInsert_Data_2_288 <= findAndInsert_Data_1_311;
                  findAndInsert_Key_3_289 <= findAndInsert_Key_2_312;
                  findAndInsert_Data_3_292 <= findAndInsert_Data_2_315;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 3;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (findAndInsert_size_301)
                0: begin
                  findAndInsert_size_274 <= findAndInsert_size_274 + 0;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                1: begin
                  findAndInsert_Key_2_285 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_2_288 <= findAndInsert_Data_0_307;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 1;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                2: begin
                  findAndInsert_Key_2_285 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_2_288 <= findAndInsert_Data_0_307;
                  findAndInsert_Key_3_289 <= findAndInsert_Key_1_308;
                  findAndInsert_Data_3_292 <= findAndInsert_Data_1_311;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 2;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (findAndInsert_size_301)
                0: begin
                  findAndInsert_size_274 <= findAndInsert_size_274 + 0;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                1: begin
                  findAndInsert_Key_3_289 <= findAndInsert_Key_0_304;
                  findAndInsert_Data_3_292 <= findAndInsert_Data_0_307;
                  findAndInsert_size_274 <= findAndInsert_size_274 + 1;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (findAndInsert_size_301)
                0: begin
                  findAndInsert_size_274 <= findAndInsert_size_274 + 0;
                  findAndInsert_MergeSuccess_299 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:1214:<init>|  Btree.java:1213:merge|  Btree.java:1902:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        375: begin
          if (findAndInsert_MergeSuccess_299 == 0) begin
            findAndInsert_pc <= 398;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0599:<init>|  Chip.java:0598:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        376: begin
          findAndInsert_size_1 <= findAndInsert_size_1-1;
          case (findAndInsert_j_48)
            0: begin
              findAndInsert_Key_39 <= findAndInsert_Key_0_4;
              findAndInsert_Data_41 <= findAndInsert_Data_0_7;
            end
            1: begin
              findAndInsert_Key_39 <= findAndInsert_Key_1_8;
              findAndInsert_Data_41 <= findAndInsert_Data_1_11;
            end
            2: begin
              findAndInsert_Key_39 <= findAndInsert_Key_2_12;
              findAndInsert_Data_41 <= findAndInsert_Data_2_15;
            end
            3: begin
              findAndInsert_Key_39 <= findAndInsert_Key_3_16;
              findAndInsert_Data_41 <= findAndInsert_Data_3_19;
            end
          endcase
          if (0>= findAndInsert_j_48) begin
            findAndInsert_Key_0_4 <= findAndInsert_Key_1_8;
            findAndInsert_Data_0_7 <= findAndInsert_Data_1_11;
          end
          if (1>= findAndInsert_j_48) begin
            findAndInsert_Key_1_8 <= findAndInsert_Key_2_12;
            findAndInsert_Data_1_11 <= findAndInsert_Data_2_15;
          end
          if (2>= findAndInsert_j_48) begin
            findAndInsert_Key_2_12 <= findAndInsert_Key_3_16;
            findAndInsert_Data_2_15 <= findAndInsert_Data_3_19;
          end
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0744:<init>|  Btree.java:0743:RemoveElementAt|  Btree.java:1906:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        377: begin
          case (findAndInsert_j_48)
            0: begin
              findAndInsert_Key_39 <= findAndInsert_Key_0_4;
              findAndInsert_Data_41 <= findAndInsert_Data_0_7;
            end
            1: begin
              findAndInsert_Key_39 <= findAndInsert_Key_1_8;
              findAndInsert_Data_41 <= findAndInsert_Data_1_11;
            end
            2: begin
              findAndInsert_Key_39 <= findAndInsert_Key_2_12;
              findAndInsert_Data_41 <= findAndInsert_Data_2_15;
            end
            3: begin
              findAndInsert_Key_39 <= findAndInsert_Key_3_16;
              findAndInsert_Data_41 <= findAndInsert_Data_3_19;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0585:<init>|  Btree.java:0584:ElementAt|  Btree.java:1907:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        378: begin
          if (findAndInsert_j_48 == findAndInsert_size_1) begin
            findAndInsert_size_1 <= findAndInsert_size_1+1;
          end
          case (findAndInsert_j_48)
            0: begin
              findAndInsert_Key_0_4 <= findAndInsert_Key_39;
              findAndInsert_Data_0_7 <= findAndInsert_indexLeft_329;
            end
            1: begin
              findAndInsert_Key_1_8 <= findAndInsert_Key_39;
              findAndInsert_Data_1_11 <= findAndInsert_indexLeft_329;
            end
            2: begin
              findAndInsert_Key_2_12 <= findAndInsert_Key_39;
              findAndInsert_Data_2_15 <= findAndInsert_indexLeft_329;
            end
            3: begin
              findAndInsert_Key_3_16 <= findAndInsert_Key_39;
              findAndInsert_Data_3_19 <= findAndInsert_indexLeft_329;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0627:<init>|  Btree.java:0626:SetElementAt|  Btree.java:1908:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        379: begin
          findAndInsert_success_332 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0795:<init>|  Chip.java:0794:One|  Btree.java:1909:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        380: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_273;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_274;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_273;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_277;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_281;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_285;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_289;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_273;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_280;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_284;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_288;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_292;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1910:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        381: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1910:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        382: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1910:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        383: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1910:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        384: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_0;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_1;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_0;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_4;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_8;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_12;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_16;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_0;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_7;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_11;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_15;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_19;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0315:<init>|  Btree.java:0314:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1911:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        385: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1911:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        386: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1911:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        387: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0333:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1911:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        388: begin
          findAndInsert_root_335 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:0788:<init>|  Chip.java:0787:Zero|  Btree.java:0128:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        389: begin
          findAndInsert_freeNext_9_index_168 <= findAndInsert_root_335;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1278:<init>|  Chip.java:1277:ExecuteTransaction|  Btree.java:0129:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        390: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1285:<init>|  Chip.java:1284:waitResultOfTransaction|  Btree.java:0130:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        391: begin
          findAndInsert_next_334 <= freeNext_freeNext_9_result_0;
          findAndInsert_freeNext_10_index_169 <= findAndInsert_root_335;
          findAndInsert_freeNext_10_value_170 <= findAndInsert_indexRight_330;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_isFree_336 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Btree.java:0133:<init>|  Btree.java:0132:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        392: begin
          findAndInsert_stuckIsFree_11_index_171 <= findAndInsert_indexRight_330;
          findAndInsert_stuckIsFree_11_value_172 <= findAndInsert_isFree_336;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1341:<init>|  Chip.java:1340:ExecuteTransaction|  Btree.java:0145:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        393: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0146:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        394: begin
          findAndInsert_freeNext_10_index_169 <= findAndInsert_indexRight_330;
          findAndInsert_freeNext_10_value_170 <= findAndInsert_next_334;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0508:<init>|  Chip.java:1341:<init>|  Chip.java:1340:ExecuteTransaction|  Btree.java:0147:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        395: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        396: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1348:<init>|  Chip.java:1347:waitResultOfTransaction|  Btree.java:0149:free|  Btree.java:1912:Then|  Chip.java:0606:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        397: begin
          findAndInsert_pc <= 398;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0608:<init>|  Chip.java:0607:<init>|  Btree.java:1905:<init>|  Btree.java:1904:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        398: begin
          findAndInsert_pc <= 399;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1901:<init>|  Btree.java:1900:Leaf|  Btree.java:1411:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        399: begin
          findAndInsert_pc <= 400;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0567:<init>|  Chip.java:0566:GOto|  Btree.java:1412:code|  Chip.java:0526:<init>|  Btree.java:1393:<init>|  Btree.java:1392:code|  Chip.java:0526:<init>|  Btree.java:1390:<init>|  Btree.java:1389:<init>|  Btree.java:1899:<init>|  Btree.java:1898:code|  Chip.java:0526:<init>|  Btree.java:1877:<init>|  Btree.java:1876:mergeLeavesNotTop|  Btree.java:4187:test_mergeLeavesNotTop|  Btree.java:7044:oldTests|  Btree.java:7064:newTests|  Btree.java:7070:main|");
            $fclose(f);
          end
        end
        default: findAndInsert_stop <= 1;
      endcase
    end
  end
  task chipPrint;
    begin
      integer o;
      o = $fopen("verilog/trace_verilog.txt", "a");
      if (!o) o = $fopen("../verilog/trace_verilog.txt", "a");
      if (!o) $display("Cannot create trace folder: verilog/trace_verilog.txt");
      $fwrite(o, "Chip: %-16s step: %1d, maxSteps: %1d, running: %1d\n", "Btree", step, maxSteps, !stop);
      $fwrite(o, "  Processes:\n");

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 0, "stuckIsLeaf", 1, stuckIsLeaf_pc, stuckIsLeaf_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsLeaf_memory[0]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[1]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[2]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[3]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[4]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[5]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[6]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[7]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[8]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[9]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[10]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[11]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[12]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[13]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[14]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[15]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[16]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[17]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[18]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[19]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[20]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[21]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[22]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[23]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[24]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[25]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[26]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[27]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[28]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[29]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[30]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckIsLeaf_7", stuckIsLeaf_7_requestedAt, stuckIsLeaf_7_finishedAt, stuckIsLeaf_stuckIsLeaf_7_returnCode, (stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step), (stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsLeaf_7_index_35", findAndInsert_stuckIsLeaf_7_index_35);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsLeaf_8", stuckIsLeaf_8_requestedAt, stuckIsLeaf_8_finishedAt, stuckIsLeaf_stuckIsLeaf_8_returnCode, (stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step), (stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsLeaf_8_index_36", findAndInsert_stuckIsLeaf_8_index_36);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsLeaf_8_value_37", findAndInsert_stuckIsLeaf_8_value_37);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 1, "stuckIsFree", 1, stuckIsFree_pc, stuckIsFree_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsFree_memory[0]);
      $fwrite(o, ", %2d", stuckIsFree_memory[1]);
      $fwrite(o, ", %2d", stuckIsFree_memory[2]);
      $fwrite(o, ", %2d", stuckIsFree_memory[3]);
      $fwrite(o, ", %2d", stuckIsFree_memory[4]);
      $fwrite(o, ", %2d", stuckIsFree_memory[5]);
      $fwrite(o, ", %2d", stuckIsFree_memory[6]);
      $fwrite(o, ", %2d", stuckIsFree_memory[7]);
      $fwrite(o, ", %2d", stuckIsFree_memory[8]);
      $fwrite(o, ", %2d", stuckIsFree_memory[9]);
      $fwrite(o, ", %2d", stuckIsFree_memory[10]);
      $fwrite(o, ", %2d", stuckIsFree_memory[11]);
      $fwrite(o, ", %2d", stuckIsFree_memory[12]);
      $fwrite(o, ", %2d", stuckIsFree_memory[13]);
      $fwrite(o, ", %2d", stuckIsFree_memory[14]);
      $fwrite(o, ", %2d", stuckIsFree_memory[15]);
      $fwrite(o, ", %2d", stuckIsFree_memory[16]);
      $fwrite(o, ", %2d", stuckIsFree_memory[17]);
      $fwrite(o, ", %2d", stuckIsFree_memory[18]);
      $fwrite(o, ", %2d", stuckIsFree_memory[19]);
      $fwrite(o, ", %2d", stuckIsFree_memory[20]);
      $fwrite(o, ", %2d", stuckIsFree_memory[21]);
      $fwrite(o, ", %2d", stuckIsFree_memory[22]);
      $fwrite(o, ", %2d", stuckIsFree_memory[23]);
      $fwrite(o, ", %2d", stuckIsFree_memory[24]);
      $fwrite(o, ", %2d", stuckIsFree_memory[25]);
      $fwrite(o, ", %2d", stuckIsFree_memory[26]);
      $fwrite(o, ", %2d", stuckIsFree_memory[27]);
      $fwrite(o, ", %2d", stuckIsFree_memory[28]);
      $fwrite(o, ", %2d", stuckIsFree_memory[29]);
      $fwrite(o, ", %2d", stuckIsFree_memory[30]);
      $fwrite(o, ", %2d", stuckIsFree_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsFree_11", stuckIsFree_11_requestedAt, stuckIsFree_11_finishedAt, stuckIsFree_stuckIsFree_11_returnCode, (stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step), (stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsFree_11_index_171", findAndInsert_stuckIsFree_11_index_171);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsFree_11_value_172", findAndInsert_stuckIsFree_11_value_172);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 2, "freeNext", 1, freeNext_pc, freeNext_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 6, 1);
      $fwrite(o, "        %2d", freeNext_memory[0]);
      $fwrite(o, ", %2d", freeNext_memory[1]);
      $fwrite(o, ", %2d", freeNext_memory[2]);
      $fwrite(o, ", %2d", freeNext_memory[3]);
      $fwrite(o, ", %2d", freeNext_memory[4]);
      $fwrite(o, ", %2d", freeNext_memory[5]);
      $fwrite(o, ", %2d", freeNext_memory[6]);
      $fwrite(o, ", %2d", freeNext_memory[7]);
      $fwrite(o, ", %2d", freeNext_memory[8]);
      $fwrite(o, ", %2d", freeNext_memory[9]);
      $fwrite(o, ", %2d", freeNext_memory[10]);
      $fwrite(o, ", %2d", freeNext_memory[11]);
      $fwrite(o, ", %2d", freeNext_memory[12]);
      $fwrite(o, ", %2d", freeNext_memory[13]);
      $fwrite(o, ", %2d", freeNext_memory[14]);
      $fwrite(o, ", %2d", freeNext_memory[15]);
      $fwrite(o, ", %2d", freeNext_memory[16]);
      $fwrite(o, ", %2d", freeNext_memory[17]);
      $fwrite(o, ", %2d", freeNext_memory[18]);
      $fwrite(o, ", %2d", freeNext_memory[19]);
      $fwrite(o, ", %2d", freeNext_memory[20]);
      $fwrite(o, ", %2d", freeNext_memory[21]);
      $fwrite(o, ", %2d", freeNext_memory[22]);
      $fwrite(o, ", %2d", freeNext_memory[23]);
      $fwrite(o, ", %2d", freeNext_memory[24]);
      $fwrite(o, ", %2d", freeNext_memory[25]);
      $fwrite(o, ", %2d", freeNext_memory[26]);
      $fwrite(o, ", %2d", freeNext_memory[27]);
      $fwrite(o, ", %2d", freeNext_memory[28]);
      $fwrite(o, ", %2d", freeNext_memory[29]);
      $fwrite(o, ", %2d", freeNext_memory[30]);
      $fwrite(o, ", %2d", freeNext_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "freeNext_9", freeNext_9_requestedAt, freeNext_9_finishedAt, freeNext_freeNext_9_returnCode, (freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step), (freeNext_9_requestedAt < freeNext_9_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_freeNext_9_index_168", findAndInsert_freeNext_9_index_168);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "freeNext_10", freeNext_10_requestedAt, freeNext_10_finishedAt, freeNext_freeNext_10_returnCode, (freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step), (freeNext_10_requestedAt < freeNext_10_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_freeNext_10_index_169", findAndInsert_freeNext_10_index_169);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_freeNext_10_value_170", findAndInsert_freeNext_10_value_170);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 3, "stuckSize", 1, stuckSize_pc, stuckSize_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 3, 1);
      $fwrite(o, "        %2d", stuckSize_memory[0]);
      $fwrite(o, ", %2d", stuckSize_memory[1]);
      $fwrite(o, ", %2d", stuckSize_memory[2]);
      $fwrite(o, ", %2d", stuckSize_memory[3]);
      $fwrite(o, ", %2d", stuckSize_memory[4]);
      $fwrite(o, ", %2d", stuckSize_memory[5]);
      $fwrite(o, ", %2d", stuckSize_memory[6]);
      $fwrite(o, ", %2d", stuckSize_memory[7]);
      $fwrite(o, ", %2d", stuckSize_memory[8]);
      $fwrite(o, ", %2d", stuckSize_memory[9]);
      $fwrite(o, ", %2d", stuckSize_memory[10]);
      $fwrite(o, ", %2d", stuckSize_memory[11]);
      $fwrite(o, ", %2d", stuckSize_memory[12]);
      $fwrite(o, ", %2d", stuckSize_memory[13]);
      $fwrite(o, ", %2d", stuckSize_memory[14]);
      $fwrite(o, ", %2d", stuckSize_memory[15]);
      $fwrite(o, ", %2d", stuckSize_memory[16]);
      $fwrite(o, ", %2d", stuckSize_memory[17]);
      $fwrite(o, ", %2d", stuckSize_memory[18]);
      $fwrite(o, ", %2d", stuckSize_memory[19]);
      $fwrite(o, ", %2d", stuckSize_memory[20]);
      $fwrite(o, ", %2d", stuckSize_memory[21]);
      $fwrite(o, ", %2d", stuckSize_memory[22]);
      $fwrite(o, ", %2d", stuckSize_memory[23]);
      $fwrite(o, ", %2d", stuckSize_memory[24]);
      $fwrite(o, ", %2d", stuckSize_memory[25]);
      $fwrite(o, ", %2d", stuckSize_memory[26]);
      $fwrite(o, ", %2d", stuckSize_memory[27]);
      $fwrite(o, ", %2d", stuckSize_memory[28]);
      $fwrite(o, ", %2d", stuckSize_memory[29]);
      $fwrite(o, ", %2d", stuckSize_memory[30]);
      $fwrite(o, ", %2d", stuckSize_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckSize_5", stuckSize_5_requestedAt, stuckSize_5_finishedAt, stuckSize_stuckSize_5_returnCode, (stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step), (stuckSize_5_requestedAt < stuckSize_5_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckSize_5_index_32", findAndInsert_stuckSize_5_index_32);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckSize_6", stuckSize_6_requestedAt, stuckSize_6_finishedAt, stuckSize_stuckSize_6_returnCode, (stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step), (stuckSize_6_requestedAt < stuckSize_6_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckSize_6_index_33", findAndInsert_stuckSize_6_index_33);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckSize_6_value_34", findAndInsert_stuckSize_6_value_34);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 4, "stuckKeys", 1, stuckKeys_pc, stuckKeys_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckKeys_memory[0]);
      $fwrite(o, ", %2d", stuckKeys_memory[1]);
      $fwrite(o, ", %2d", stuckKeys_memory[2]);
      $fwrite(o, ", %2d", stuckKeys_memory[3]);
      $fwrite(o, ", %2d", stuckKeys_memory[4]);
      $fwrite(o, ", %2d", stuckKeys_memory[5]);
      $fwrite(o, ", %2d", stuckKeys_memory[6]);
      $fwrite(o, ", %2d", stuckKeys_memory[7]);
      $fwrite(o, ", %2d", stuckKeys_memory[8]);
      $fwrite(o, ", %2d", stuckKeys_memory[9]);
      $fwrite(o, ", %2d", stuckKeys_memory[10]);
      $fwrite(o, ", %2d", stuckKeys_memory[11]);
      $fwrite(o, ", %2d", stuckKeys_memory[12]);
      $fwrite(o, ", %2d", stuckKeys_memory[13]);
      $fwrite(o, ", %2d", stuckKeys_memory[14]);
      $fwrite(o, ", %2d", stuckKeys_memory[15]);
      $fwrite(o, ", %2d", stuckKeys_memory[16]);
      $fwrite(o, ", %2d", stuckKeys_memory[17]);
      $fwrite(o, ", %2d", stuckKeys_memory[18]);
      $fwrite(o, ", %2d", stuckKeys_memory[19]);
      $fwrite(o, ", %2d", stuckKeys_memory[20]);
      $fwrite(o, ", %2d", stuckKeys_memory[21]);
      $fwrite(o, ", %2d", stuckKeys_memory[22]);
      $fwrite(o, ", %2d", stuckKeys_memory[23]);
      $fwrite(o, ", %2d", stuckKeys_memory[24]);
      $fwrite(o, ", %2d", stuckKeys_memory[25]);
      $fwrite(o, ", %2d", stuckKeys_memory[26]);
      $fwrite(o, ", %2d", stuckKeys_memory[27]);
      $fwrite(o, ", %2d", stuckKeys_memory[28]);
      $fwrite(o, ", %2d", stuckKeys_memory[29]);
      $fwrite(o, ", %2d", stuckKeys_memory[30]);
      $fwrite(o, ", %2d", stuckKeys_memory[31]);
      $fwrite(o, ", %2d", stuckKeys_memory[32]);
      $fwrite(o, ", %2d", stuckKeys_memory[33]);
      $fwrite(o, ", %2d", stuckKeys_memory[34]);
      $fwrite(o, ", %2d", stuckKeys_memory[35]);
      $fwrite(o, ", %2d", stuckKeys_memory[36]);
      $fwrite(o, ", %2d", stuckKeys_memory[37]);
      $fwrite(o, ", %2d", stuckKeys_memory[38]);
      $fwrite(o, ", %2d", stuckKeys_memory[39]);
      $fwrite(o, ", %2d", stuckKeys_memory[40]);
      $fwrite(o, ", %2d", stuckKeys_memory[41]);
      $fwrite(o, ", %2d", stuckKeys_memory[42]);
      $fwrite(o, ", %2d", stuckKeys_memory[43]);
      $fwrite(o, ", %2d", stuckKeys_memory[44]);
      $fwrite(o, ", %2d", stuckKeys_memory[45]);
      $fwrite(o, ", %2d", stuckKeys_memory[46]);
      $fwrite(o, ", %2d", stuckKeys_memory[47]);
      $fwrite(o, ", %2d", stuckKeys_memory[48]);
      $fwrite(o, ", %2d", stuckKeys_memory[49]);
      $fwrite(o, ", %2d", stuckKeys_memory[50]);
      $fwrite(o, ", %2d", stuckKeys_memory[51]);
      $fwrite(o, ", %2d", stuckKeys_memory[52]);
      $fwrite(o, ", %2d", stuckKeys_memory[53]);
      $fwrite(o, ", %2d", stuckKeys_memory[54]);
      $fwrite(o, ", %2d", stuckKeys_memory[55]);
      $fwrite(o, ", %2d", stuckKeys_memory[56]);
      $fwrite(o, ", %2d", stuckKeys_memory[57]);
      $fwrite(o, ", %2d", stuckKeys_memory[58]);
      $fwrite(o, ", %2d", stuckKeys_memory[59]);
      $fwrite(o, ", %2d", stuckKeys_memory[60]);
      $fwrite(o, ", %2d", stuckKeys_memory[61]);
      $fwrite(o, ", %2d", stuckKeys_memory[62]);
      $fwrite(o, ", %2d", stuckKeys_memory[63]);
      $fwrite(o, ", %2d", stuckKeys_memory[64]);
      $fwrite(o, ", %2d", stuckKeys_memory[65]);
      $fwrite(o, ", %2d", stuckKeys_memory[66]);
      $fwrite(o, ", %2d", stuckKeys_memory[67]);
      $fwrite(o, ", %2d", stuckKeys_memory[68]);
      $fwrite(o, ", %2d", stuckKeys_memory[69]);
      $fwrite(o, ", %2d", stuckKeys_memory[70]);
      $fwrite(o, ", %2d", stuckKeys_memory[71]);
      $fwrite(o, ", %2d", stuckKeys_memory[72]);
      $fwrite(o, ", %2d", stuckKeys_memory[73]);
      $fwrite(o, ", %2d", stuckKeys_memory[74]);
      $fwrite(o, ", %2d", stuckKeys_memory[75]);
      $fwrite(o, ", %2d", stuckKeys_memory[76]);
      $fwrite(o, ", %2d", stuckKeys_memory[77]);
      $fwrite(o, ", %2d", stuckKeys_memory[78]);
      $fwrite(o, ", %2d", stuckKeys_memory[79]);
      $fwrite(o, ", %2d", stuckKeys_memory[80]);
      $fwrite(o, ", %2d", stuckKeys_memory[81]);
      $fwrite(o, ", %2d", stuckKeys_memory[82]);
      $fwrite(o, ", %2d", stuckKeys_memory[83]);
      $fwrite(o, ", %2d", stuckKeys_memory[84]);
      $fwrite(o, ", %2d", stuckKeys_memory[85]);
      $fwrite(o, ", %2d", stuckKeys_memory[86]);
      $fwrite(o, ", %2d", stuckKeys_memory[87]);
      $fwrite(o, ", %2d", stuckKeys_memory[88]);
      $fwrite(o, ", %2d", stuckKeys_memory[89]);
      $fwrite(o, ", %2d", stuckKeys_memory[90]);
      $fwrite(o, ", %2d", stuckKeys_memory[91]);
      $fwrite(o, ", %2d", stuckKeys_memory[92]);
      $fwrite(o, ", %2d", stuckKeys_memory[93]);
      $fwrite(o, ", %2d", stuckKeys_memory[94]);
      $fwrite(o, ", %2d", stuckKeys_memory[95]);
      $fwrite(o, ", %2d", stuckKeys_memory[96]);
      $fwrite(o, ", %2d", stuckKeys_memory[97]);
      $fwrite(o, ", %2d", stuckKeys_memory[98]);
      $fwrite(o, ", %2d", stuckKeys_memory[99]);
      $fwrite(o, ", %2d", stuckKeys_memory[100]);
      $fwrite(o, ", %2d", stuckKeys_memory[101]);
      $fwrite(o, ", %2d", stuckKeys_memory[102]);
      $fwrite(o, ", %2d", stuckKeys_memory[103]);
      $fwrite(o, ", %2d", stuckKeys_memory[104]);
      $fwrite(o, ", %2d", stuckKeys_memory[105]);
      $fwrite(o, ", %2d", stuckKeys_memory[106]);
      $fwrite(o, ", %2d", stuckKeys_memory[107]);
      $fwrite(o, ", %2d", stuckKeys_memory[108]);
      $fwrite(o, ", %2d", stuckKeys_memory[109]);
      $fwrite(o, ", %2d", stuckKeys_memory[110]);
      $fwrite(o, ", %2d", stuckKeys_memory[111]);
      $fwrite(o, ", %2d", stuckKeys_memory[112]);
      $fwrite(o, ", %2d", stuckKeys_memory[113]);
      $fwrite(o, ", %2d", stuckKeys_memory[114]);
      $fwrite(o, ", %2d", stuckKeys_memory[115]);
      $fwrite(o, ", %2d", stuckKeys_memory[116]);
      $fwrite(o, ", %2d", stuckKeys_memory[117]);
      $fwrite(o, ", %2d", stuckKeys_memory[118]);
      $fwrite(o, ", %2d", stuckKeys_memory[119]);
      $fwrite(o, ", %2d", stuckKeys_memory[120]);
      $fwrite(o, ", %2d", stuckKeys_memory[121]);
      $fwrite(o, ", %2d", stuckKeys_memory[122]);
      $fwrite(o, ", %2d", stuckKeys_memory[123]);
      $fwrite(o, ", %2d", stuckKeys_memory[124]);
      $fwrite(o, ", %2d", stuckKeys_memory[125]);
      $fwrite(o, ", %2d", stuckKeys_memory[126]);
      $fwrite(o, ", %2d", stuckKeys_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckKeys_1", stuckKeys_1_requestedAt, stuckKeys_1_finishedAt, stuckKeys_stuckKeys_1_returnCode, (stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step), (stuckKeys_1_requestedAt < stuckKeys_1_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_1_index_20", findAndInsert_stuckKeys_1_index_20);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckKeys_2", stuckKeys_2_requestedAt, stuckKeys_2_finishedAt, stuckKeys_stuckKeys_2_returnCode, (stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step), (stuckKeys_2_requestedAt < stuckKeys_2_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_index_21", findAndInsert_stuckKeys_2_index_21);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_22", findAndInsert_stuckKeys_2_value_22);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_23", findAndInsert_stuckKeys_2_value_23);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_24", findAndInsert_stuckKeys_2_value_24);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_25", findAndInsert_stuckKeys_2_value_25);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 5, "stuckData", 1, stuckData_pc, stuckData_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckData_memory[0]);
      $fwrite(o, ", %2d", stuckData_memory[1]);
      $fwrite(o, ", %2d", stuckData_memory[2]);
      $fwrite(o, ", %2d", stuckData_memory[3]);
      $fwrite(o, ", %2d", stuckData_memory[4]);
      $fwrite(o, ", %2d", stuckData_memory[5]);
      $fwrite(o, ", %2d", stuckData_memory[6]);
      $fwrite(o, ", %2d", stuckData_memory[7]);
      $fwrite(o, ", %2d", stuckData_memory[8]);
      $fwrite(o, ", %2d", stuckData_memory[9]);
      $fwrite(o, ", %2d", stuckData_memory[10]);
      $fwrite(o, ", %2d", stuckData_memory[11]);
      $fwrite(o, ", %2d", stuckData_memory[12]);
      $fwrite(o, ", %2d", stuckData_memory[13]);
      $fwrite(o, ", %2d", stuckData_memory[14]);
      $fwrite(o, ", %2d", stuckData_memory[15]);
      $fwrite(o, ", %2d", stuckData_memory[16]);
      $fwrite(o, ", %2d", stuckData_memory[17]);
      $fwrite(o, ", %2d", stuckData_memory[18]);
      $fwrite(o, ", %2d", stuckData_memory[19]);
      $fwrite(o, ", %2d", stuckData_memory[20]);
      $fwrite(o, ", %2d", stuckData_memory[21]);
      $fwrite(o, ", %2d", stuckData_memory[22]);
      $fwrite(o, ", %2d", stuckData_memory[23]);
      $fwrite(o, ", %2d", stuckData_memory[24]);
      $fwrite(o, ", %2d", stuckData_memory[25]);
      $fwrite(o, ", %2d", stuckData_memory[26]);
      $fwrite(o, ", %2d", stuckData_memory[27]);
      $fwrite(o, ", %2d", stuckData_memory[28]);
      $fwrite(o, ", %2d", stuckData_memory[29]);
      $fwrite(o, ", %2d", stuckData_memory[30]);
      $fwrite(o, ", %2d", stuckData_memory[31]);
      $fwrite(o, ", %2d", stuckData_memory[32]);
      $fwrite(o, ", %2d", stuckData_memory[33]);
      $fwrite(o, ", %2d", stuckData_memory[34]);
      $fwrite(o, ", %2d", stuckData_memory[35]);
      $fwrite(o, ", %2d", stuckData_memory[36]);
      $fwrite(o, ", %2d", stuckData_memory[37]);
      $fwrite(o, ", %2d", stuckData_memory[38]);
      $fwrite(o, ", %2d", stuckData_memory[39]);
      $fwrite(o, ", %2d", stuckData_memory[40]);
      $fwrite(o, ", %2d", stuckData_memory[41]);
      $fwrite(o, ", %2d", stuckData_memory[42]);
      $fwrite(o, ", %2d", stuckData_memory[43]);
      $fwrite(o, ", %2d", stuckData_memory[44]);
      $fwrite(o, ", %2d", stuckData_memory[45]);
      $fwrite(o, ", %2d", stuckData_memory[46]);
      $fwrite(o, ", %2d", stuckData_memory[47]);
      $fwrite(o, ", %2d", stuckData_memory[48]);
      $fwrite(o, ", %2d", stuckData_memory[49]);
      $fwrite(o, ", %2d", stuckData_memory[50]);
      $fwrite(o, ", %2d", stuckData_memory[51]);
      $fwrite(o, ", %2d", stuckData_memory[52]);
      $fwrite(o, ", %2d", stuckData_memory[53]);
      $fwrite(o, ", %2d", stuckData_memory[54]);
      $fwrite(o, ", %2d", stuckData_memory[55]);
      $fwrite(o, ", %2d", stuckData_memory[56]);
      $fwrite(o, ", %2d", stuckData_memory[57]);
      $fwrite(o, ", %2d", stuckData_memory[58]);
      $fwrite(o, ", %2d", stuckData_memory[59]);
      $fwrite(o, ", %2d", stuckData_memory[60]);
      $fwrite(o, ", %2d", stuckData_memory[61]);
      $fwrite(o, ", %2d", stuckData_memory[62]);
      $fwrite(o, ", %2d", stuckData_memory[63]);
      $fwrite(o, ", %2d", stuckData_memory[64]);
      $fwrite(o, ", %2d", stuckData_memory[65]);
      $fwrite(o, ", %2d", stuckData_memory[66]);
      $fwrite(o, ", %2d", stuckData_memory[67]);
      $fwrite(o, ", %2d", stuckData_memory[68]);
      $fwrite(o, ", %2d", stuckData_memory[69]);
      $fwrite(o, ", %2d", stuckData_memory[70]);
      $fwrite(o, ", %2d", stuckData_memory[71]);
      $fwrite(o, ", %2d", stuckData_memory[72]);
      $fwrite(o, ", %2d", stuckData_memory[73]);
      $fwrite(o, ", %2d", stuckData_memory[74]);
      $fwrite(o, ", %2d", stuckData_memory[75]);
      $fwrite(o, ", %2d", stuckData_memory[76]);
      $fwrite(o, ", %2d", stuckData_memory[77]);
      $fwrite(o, ", %2d", stuckData_memory[78]);
      $fwrite(o, ", %2d", stuckData_memory[79]);
      $fwrite(o, ", %2d", stuckData_memory[80]);
      $fwrite(o, ", %2d", stuckData_memory[81]);
      $fwrite(o, ", %2d", stuckData_memory[82]);
      $fwrite(o, ", %2d", stuckData_memory[83]);
      $fwrite(o, ", %2d", stuckData_memory[84]);
      $fwrite(o, ", %2d", stuckData_memory[85]);
      $fwrite(o, ", %2d", stuckData_memory[86]);
      $fwrite(o, ", %2d", stuckData_memory[87]);
      $fwrite(o, ", %2d", stuckData_memory[88]);
      $fwrite(o, ", %2d", stuckData_memory[89]);
      $fwrite(o, ", %2d", stuckData_memory[90]);
      $fwrite(o, ", %2d", stuckData_memory[91]);
      $fwrite(o, ", %2d", stuckData_memory[92]);
      $fwrite(o, ", %2d", stuckData_memory[93]);
      $fwrite(o, ", %2d", stuckData_memory[94]);
      $fwrite(o, ", %2d", stuckData_memory[95]);
      $fwrite(o, ", %2d", stuckData_memory[96]);
      $fwrite(o, ", %2d", stuckData_memory[97]);
      $fwrite(o, ", %2d", stuckData_memory[98]);
      $fwrite(o, ", %2d", stuckData_memory[99]);
      $fwrite(o, ", %2d", stuckData_memory[100]);
      $fwrite(o, ", %2d", stuckData_memory[101]);
      $fwrite(o, ", %2d", stuckData_memory[102]);
      $fwrite(o, ", %2d", stuckData_memory[103]);
      $fwrite(o, ", %2d", stuckData_memory[104]);
      $fwrite(o, ", %2d", stuckData_memory[105]);
      $fwrite(o, ", %2d", stuckData_memory[106]);
      $fwrite(o, ", %2d", stuckData_memory[107]);
      $fwrite(o, ", %2d", stuckData_memory[108]);
      $fwrite(o, ", %2d", stuckData_memory[109]);
      $fwrite(o, ", %2d", stuckData_memory[110]);
      $fwrite(o, ", %2d", stuckData_memory[111]);
      $fwrite(o, ", %2d", stuckData_memory[112]);
      $fwrite(o, ", %2d", stuckData_memory[113]);
      $fwrite(o, ", %2d", stuckData_memory[114]);
      $fwrite(o, ", %2d", stuckData_memory[115]);
      $fwrite(o, ", %2d", stuckData_memory[116]);
      $fwrite(o, ", %2d", stuckData_memory[117]);
      $fwrite(o, ", %2d", stuckData_memory[118]);
      $fwrite(o, ", %2d", stuckData_memory[119]);
      $fwrite(o, ", %2d", stuckData_memory[120]);
      $fwrite(o, ", %2d", stuckData_memory[121]);
      $fwrite(o, ", %2d", stuckData_memory[122]);
      $fwrite(o, ", %2d", stuckData_memory[123]);
      $fwrite(o, ", %2d", stuckData_memory[124]);
      $fwrite(o, ", %2d", stuckData_memory[125]);
      $fwrite(o, ", %2d", stuckData_memory[126]);
      $fwrite(o, ", %2d", stuckData_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckData_3", stuckData_3_requestedAt, stuckData_3_finishedAt, stuckData_stuckData_3_returnCode, (stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step), (stuckData_3_requestedAt < stuckData_3_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_3_index_26", findAndInsert_stuckData_3_index_26);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckData_4", stuckData_4_requestedAt, stuckData_4_finishedAt, stuckData_stuckData_4_returnCode, (stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step), (stuckData_4_requestedAt < stuckData_4_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_index_27", findAndInsert_stuckData_4_index_27);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_28", findAndInsert_stuckData_4_value_28);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_29", findAndInsert_stuckData_4_value_29);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_30", findAndInsert_stuckData_4_value_30);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_31", findAndInsert_stuckData_4_value_31);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 6, "findAndInsert", 400, findAndInsert_pc, findAndInsert_returnCode);
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_0", findAndInsert_index_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_1", findAndInsert_size_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_2", findAndInsert_isLeaf_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_3", findAndInsert_nextFree_3);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_4", findAndInsert_Key_0_4);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_5", findAndInsert_KeyCompares_0_5);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_6", findAndInsert_KeyCollapse_0_6);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_7", findAndInsert_Data_0_7);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_8", findAndInsert_Key_1_8);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_9", findAndInsert_KeyCompares_1_9);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_10", findAndInsert_KeyCollapse_1_10);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_11", findAndInsert_Data_1_11);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_12", findAndInsert_Key_2_12);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_13", findAndInsert_KeyCompares_2_13);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_14", findAndInsert_KeyCollapse_2_14);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_15", findAndInsert_Data_2_15);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_16", findAndInsert_Key_3_16);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_17", findAndInsert_KeyCompares_3_17);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_18", findAndInsert_KeyCollapse_3_18);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_19", findAndInsert_Data_3_19);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_1_index_20", findAndInsert_stuckKeys_1_index_20);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_index_21", findAndInsert_stuckKeys_2_index_21);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_22", findAndInsert_stuckKeys_2_value_22);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_23", findAndInsert_stuckKeys_2_value_23);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_24", findAndInsert_stuckKeys_2_value_24);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_25", findAndInsert_stuckKeys_2_value_25);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_3_index_26", findAndInsert_stuckData_3_index_26);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_index_27", findAndInsert_stuckData_4_index_27);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_28", findAndInsert_stuckData_4_value_28);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_29", findAndInsert_stuckData_4_value_29);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_30", findAndInsert_stuckData_4_value_30);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_31", findAndInsert_stuckData_4_value_31);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckSize_5_index_32", findAndInsert_stuckSize_5_index_32);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckSize_6_index_33", findAndInsert_stuckSize_6_index_33);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckSize_6_value_34", findAndInsert_stuckSize_6_value_34);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsLeaf_7_index_35", findAndInsert_stuckIsLeaf_7_index_35);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsLeaf_8_index_36", findAndInsert_stuckIsLeaf_8_index_36);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsLeaf_8_value_37", findAndInsert_stuckIsLeaf_8_value_37);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_38", findAndInsert_Found_38);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_39", findAndInsert_Key_39);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_40", findAndInsert_FoundKey_40);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_41", findAndInsert_Data_41);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_42", findAndInsert_BtreeIndex_42);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_43", findAndInsert_StuckIndex_43);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_44", findAndInsert_MergeSuccess_44);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_k_45", findAndInsert_k_45);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_d_46", findAndInsert_d_46);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_47", findAndInsert_i_47);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_j_48", findAndInsert_j_48);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_49", findAndInsert_index_49);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_50", findAndInsert_size_50);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_51", findAndInsert_isLeaf_51);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_52", findAndInsert_nextFree_52);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_53", findAndInsert_Key_0_53);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_54", findAndInsert_KeyCompares_0_54);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_55", findAndInsert_KeyCollapse_0_55);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_56", findAndInsert_Data_0_56);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_57", findAndInsert_Key_1_57);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_58", findAndInsert_KeyCompares_1_58);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_59", findAndInsert_KeyCollapse_1_59);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_60", findAndInsert_Data_1_60);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_61", findAndInsert_Key_2_61);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_62", findAndInsert_KeyCompares_2_62);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_63", findAndInsert_KeyCollapse_2_63);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_64", findAndInsert_Data_2_64);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_65", findAndInsert_Key_3_65);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_66", findAndInsert_KeyCompares_3_66);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_67", findAndInsert_KeyCollapse_3_67);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_68", findAndInsert_Data_3_68);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_69", findAndInsert_Found_69);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_70", findAndInsert_Key_70);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_71", findAndInsert_FoundKey_71);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_72", findAndInsert_Data_72);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_73", findAndInsert_BtreeIndex_73);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_74", findAndInsert_StuckIndex_74);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_75", findAndInsert_MergeSuccess_75);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_76", findAndInsert_i_76);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_notFull_77", findAndInsert_notFull_77);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_78", findAndInsert_i_78);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_notFull_79", findAndInsert_notFull_79);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_80", findAndInsert_i_80);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_notFull_81", findAndInsert_notFull_81);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_82", findAndInsert_i_82);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_notFull_83", findAndInsert_notFull_83);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_84", findAndInsert_index_84);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_85", findAndInsert_size_85);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_86", findAndInsert_isLeaf_86);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_87", findAndInsert_nextFree_87);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_88", findAndInsert_Key_0_88);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_89", findAndInsert_KeyCompares_0_89);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_90", findAndInsert_KeyCollapse_0_90);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_91", findAndInsert_Data_0_91);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_92", findAndInsert_Key_1_92);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_93", findAndInsert_KeyCompares_1_93);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_94", findAndInsert_KeyCollapse_1_94);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_95", findAndInsert_Data_1_95);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_96", findAndInsert_Key_2_96);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_97", findAndInsert_KeyCompares_2_97);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_98", findAndInsert_KeyCollapse_2_98);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_99", findAndInsert_Data_2_99);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_100", findAndInsert_Key_3_100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_101", findAndInsert_KeyCompares_3_101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_102", findAndInsert_KeyCollapse_3_102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_103", findAndInsert_Data_3_103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_104", findAndInsert_Found_104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_105", findAndInsert_Key_105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_106", findAndInsert_FoundKey_106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_107", findAndInsert_Data_107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_108", findAndInsert_BtreeIndex_108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_109", findAndInsert_StuckIndex_109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_110", findAndInsert_MergeSuccess_110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_111", findAndInsert_index_111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_112", findAndInsert_size_112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_113", findAndInsert_isLeaf_113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_114", findAndInsert_nextFree_114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_115", findAndInsert_Key_0_115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_116", findAndInsert_KeyCompares_0_116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_117", findAndInsert_KeyCollapse_0_117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_118", findAndInsert_Data_0_118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_119", findAndInsert_Key_1_119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_120", findAndInsert_KeyCompares_1_120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_121", findAndInsert_KeyCollapse_1_121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_122", findAndInsert_Data_1_122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_123", findAndInsert_Key_2_123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_124", findAndInsert_KeyCompares_2_124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_125", findAndInsert_KeyCollapse_2_125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_126", findAndInsert_Data_2_126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_127", findAndInsert_Key_3_127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_128", findAndInsert_KeyCompares_3_128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_129", findAndInsert_KeyCollapse_3_129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_130", findAndInsert_Data_3_130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_131", findAndInsert_Found_131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_132", findAndInsert_Key_132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_133", findAndInsert_FoundKey_133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_134", findAndInsert_Data_134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_135", findAndInsert_BtreeIndex_135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_136", findAndInsert_StuckIndex_136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_137", findAndInsert_MergeSuccess_137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_138", findAndInsert_index_138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_139", findAndInsert_size_139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_140", findAndInsert_isLeaf_140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_141", findAndInsert_nextFree_141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_142", findAndInsert_Key_0_142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_143", findAndInsert_KeyCompares_0_143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_144", findAndInsert_KeyCollapse_0_144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_145", findAndInsert_Data_0_145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_146", findAndInsert_Key_1_146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_147", findAndInsert_KeyCompares_1_147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_148", findAndInsert_KeyCollapse_1_148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_149", findAndInsert_Data_1_149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_150", findAndInsert_Key_2_150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_151", findAndInsert_KeyCompares_2_151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_152", findAndInsert_KeyCollapse_2_152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_153", findAndInsert_Data_2_153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_154", findAndInsert_Key_3_154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_155", findAndInsert_KeyCompares_3_155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_156", findAndInsert_KeyCollapse_3_156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_157", findAndInsert_Data_3_157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_158", findAndInsert_Found_158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_159", findAndInsert_Key_159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_160", findAndInsert_FoundKey_160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_161", findAndInsert_Data_161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_162", findAndInsert_BtreeIndex_162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_163", findAndInsert_StuckIndex_163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_164", findAndInsert_MergeSuccess_164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexLeft_165", findAndInsert_indexLeft_165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexRight_166", findAndInsert_indexRight_166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_midKey_167", findAndInsert_midKey_167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_freeNext_9_index_168", findAndInsert_freeNext_9_index_168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_freeNext_10_index_169", findAndInsert_freeNext_10_index_169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_freeNext_10_value_170", findAndInsert_freeNext_10_value_170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsFree_11_index_171", findAndInsert_stuckIsFree_11_index_171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsFree_11_value_172", findAndInsert_stuckIsFree_11_value_172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_root_173", findAndInsert_root_173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_next_174", findAndInsert_next_174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_175", findAndInsert_isLeaf_175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isFree_176", findAndInsert_isFree_176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_root_177", findAndInsert_root_177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_next_178", findAndInsert_next_178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_179", findAndInsert_isLeaf_179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isFree_180", findAndInsert_isFree_180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_181", findAndInsert_i_181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_notFull_182", findAndInsert_notFull_182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_183", findAndInsert_i_183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_notFull_184", findAndInsert_notFull_184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_185", findAndInsert_index_185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_186", findAndInsert_size_186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_187", findAndInsert_isLeaf_187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_188", findAndInsert_nextFree_188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_189", findAndInsert_Key_0_189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_190", findAndInsert_KeyCompares_0_190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_191", findAndInsert_KeyCollapse_0_191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_192", findAndInsert_Data_0_192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_193", findAndInsert_Key_1_193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_194", findAndInsert_KeyCompares_1_194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_195", findAndInsert_KeyCollapse_1_195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_196", findAndInsert_Data_1_196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_197", findAndInsert_Key_2_197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_198", findAndInsert_KeyCompares_2_198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_199", findAndInsert_KeyCollapse_2_199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_200", findAndInsert_Data_2_200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_201", findAndInsert_Key_3_201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_202", findAndInsert_KeyCompares_3_202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_203", findAndInsert_KeyCollapse_3_203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_204", findAndInsert_Data_3_204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_205", findAndInsert_Found_205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_206", findAndInsert_Key_206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_207", findAndInsert_FoundKey_207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_208", findAndInsert_Data_208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_209", findAndInsert_BtreeIndex_209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_210", findAndInsert_StuckIndex_210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_211", findAndInsert_MergeSuccess_211);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_212", findAndInsert_index_212);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_213", findAndInsert_size_213);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_214", findAndInsert_isLeaf_214);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_215", findAndInsert_nextFree_215);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_216", findAndInsert_Key_0_216);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_217", findAndInsert_KeyCompares_0_217);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_218", findAndInsert_KeyCollapse_0_218);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_219", findAndInsert_Data_0_219);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_220", findAndInsert_Key_1_220);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_221", findAndInsert_KeyCompares_1_221);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_222", findAndInsert_KeyCollapse_1_222);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_223", findAndInsert_Data_1_223);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_224", findAndInsert_Key_2_224);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_225", findAndInsert_KeyCompares_2_225);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_226", findAndInsert_KeyCollapse_2_226);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_227", findAndInsert_Data_2_227);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_228", findAndInsert_Key_3_228);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_229", findAndInsert_KeyCompares_3_229);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_230", findAndInsert_KeyCollapse_3_230);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_231", findAndInsert_Data_3_231);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_232", findAndInsert_Found_232);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_233", findAndInsert_Key_233);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_234", findAndInsert_FoundKey_234);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_235", findAndInsert_Data_235);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_236", findAndInsert_BtreeIndex_236);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_237", findAndInsert_StuckIndex_237);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_238", findAndInsert_MergeSuccess_238);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_239", findAndInsert_index_239);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_240", findAndInsert_size_240);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_241", findAndInsert_isLeaf_241);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_242", findAndInsert_nextFree_242);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_243", findAndInsert_Key_0_243);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_244", findAndInsert_KeyCompares_0_244);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_245", findAndInsert_KeyCollapse_0_245);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_246", findAndInsert_Data_0_246);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_247", findAndInsert_Key_1_247);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_248", findAndInsert_KeyCompares_1_248);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_249", findAndInsert_KeyCollapse_1_249);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_250", findAndInsert_Data_1_250);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_251", findAndInsert_Key_2_251);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_252", findAndInsert_KeyCompares_2_252);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_253", findAndInsert_KeyCollapse_2_253);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_254", findAndInsert_Data_2_254);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_255", findAndInsert_Key_3_255);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_256", findAndInsert_KeyCompares_3_256);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_257", findAndInsert_KeyCollapse_3_257);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_258", findAndInsert_Data_3_258);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_259", findAndInsert_Found_259);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_260", findAndInsert_Key_260);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_261", findAndInsert_FoundKey_261);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_262", findAndInsert_Data_262);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_263", findAndInsert_BtreeIndex_263);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_264", findAndInsert_StuckIndex_264);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_265", findAndInsert_MergeSuccess_265);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childIndex_266", findAndInsert_childIndex_266);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_leftIndex_267", findAndInsert_leftIndex_267);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_midKey_268", findAndInsert_midKey_268);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_root_269", findAndInsert_root_269);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_next_270", findAndInsert_next_270);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_271", findAndInsert_isLeaf_271);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isFree_272", findAndInsert_isFree_272);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_273", findAndInsert_index_273);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_274", findAndInsert_size_274);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_275", findAndInsert_isLeaf_275);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_276", findAndInsert_nextFree_276);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_277", findAndInsert_Key_0_277);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_278", findAndInsert_KeyCompares_0_278);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_279", findAndInsert_KeyCollapse_0_279);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_280", findAndInsert_Data_0_280);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_281", findAndInsert_Key_1_281);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_282", findAndInsert_KeyCompares_1_282);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_283", findAndInsert_KeyCollapse_1_283);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_284", findAndInsert_Data_1_284);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_285", findAndInsert_Key_2_285);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_286", findAndInsert_KeyCompares_2_286);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_287", findAndInsert_KeyCollapse_2_287);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_288", findAndInsert_Data_2_288);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_289", findAndInsert_Key_3_289);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_290", findAndInsert_KeyCompares_3_290);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_291", findAndInsert_KeyCollapse_3_291);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_292", findAndInsert_Data_3_292);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_293", findAndInsert_Found_293);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_294", findAndInsert_Key_294);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_295", findAndInsert_FoundKey_295);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_296", findAndInsert_Data_296);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_297", findAndInsert_BtreeIndex_297);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_298", findAndInsert_StuckIndex_298);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_299", findAndInsert_MergeSuccess_299);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_300", findAndInsert_index_300);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_301", findAndInsert_size_301);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_302", findAndInsert_isLeaf_302);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_303", findAndInsert_nextFree_303);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_304", findAndInsert_Key_0_304);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_305", findAndInsert_KeyCompares_0_305);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_306", findAndInsert_KeyCollapse_0_306);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_307", findAndInsert_Data_0_307);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_308", findAndInsert_Key_1_308);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_309", findAndInsert_KeyCompares_1_309);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_310", findAndInsert_KeyCollapse_1_310);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_311", findAndInsert_Data_1_311);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_312", findAndInsert_Key_2_312);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_313", findAndInsert_KeyCompares_2_313);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_314", findAndInsert_KeyCollapse_2_314);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_315", findAndInsert_Data_2_315);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_316", findAndInsert_Key_3_316);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_317", findAndInsert_KeyCompares_3_317);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_318", findAndInsert_KeyCollapse_3_318);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_319", findAndInsert_Data_3_319);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_320", findAndInsert_Found_320);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_321", findAndInsert_Key_321);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_322", findAndInsert_FoundKey_322);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_323", findAndInsert_Data_323);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_324", findAndInsert_BtreeIndex_324);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_325", findAndInsert_StuckIndex_325);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_326", findAndInsert_MergeSuccess_326);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childKey_327", findAndInsert_childKey_327);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childData_328", findAndInsert_childData_328);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexLeft_329", findAndInsert_indexLeft_329);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexRight_330", findAndInsert_indexRight_330);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_midKey_331", findAndInsert_midKey_331);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_success_332", findAndInsert_success_332);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_test_333", findAndInsert_test_333);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_next_334", findAndInsert_next_334);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_root_335", findAndInsert_root_335);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isFree_336", findAndInsert_isFree_336);
      $fclose(o);
    end
  endtask
endmodule
