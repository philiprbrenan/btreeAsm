//-----------------------------------------------------------------------------
// Database on a chip test bench
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree;                                                                      // Test bench for database on a chip
  reg                    stop;                                                  // Program has stopped when this goes high
  reg                   clock;                                                  // Clock
  integer                step;                                                  // Step of the simulation
  integer            maxSteps;                                                  // Maximum number of steps to execute
  integer          returnCode;                                                  // Return code
  integer      processCurrent;                                                  // To ensure we get the same results in Java and Verilog we have to run the processes single threaded in a constant order

  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_stop||stuckData_stop||delete_stop;                                                             // Or of process stop fields

  initial begin
    returnCode = 0;
    maxSteps = 40000;
    for(step = -1; step < 0 || step < maxSteps && !stop; step = step + 1) begin // Steps below zero are run unconditionally to initialize each process so that Java and Verilog start in sync at step zero

      processCurrent = 0; clock = 0; #1; clock = 1; #1; // process_stuckIsLeaf_0000
      processCurrent = 1; clock = 0; #1; clock = 1; #1; // process_stuckIsFree_0001
      processCurrent = 2; clock = 0; #1; clock = 1; #1; // process_freeNext_0002
      processCurrent = 3; clock = 0; #1; clock = 1; #1; // process_stuckSize_0003
      processCurrent = 4; clock = 0; #1; clock = 1; #1; // process_stuckKeys_0004
      processCurrent = 5; clock = 0; #1; clock = 1; #1; // process_stuckData_0005
      processCurrent = 6; clock = 0; #1; clock = 1; #1; // process_delete_0006
      if (step >= 0) chipPrint();                                            // Steps prior to zero are for initialization to make Java and Verilog match
    end
    if (!stop) $finish(1); else $finish(0);                                // Set return code depending on whether the simulation halted
  end
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[32*1];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_7_result_0;
  integer stuckIsLeaf_7_requestedAt;
  integer stuckIsLeaf_7_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_7_returnCode;
  integer stuckIsLeaf_8_requestedAt;
  integer stuckIsLeaf_8_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_8_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  integer stuckIsLeaf_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_7_result_0 <= 0;
      stuckIsLeaf_7_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_7_returnCode <= 0;
      stuckIsLeaf_8_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_8_returnCode <= 0;
      for(stuckIsLeaf_memory_index = 0; stuckIsLeaf_memory_index < 1; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
      stuckIsLeaf_memory[1] <= 1;
      stuckIsLeaf_memory[2] <= 1;
      stuckIsLeaf_memory[3] <= 1;
      stuckIsLeaf_memory[4] <= 1;
      for(stuckIsLeaf_memory_index = 5; stuckIsLeaf_memory_index < 7; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
      stuckIsLeaf_memory[7] <= 1;
      stuckIsLeaf_memory[8] <= 1;
      stuckIsLeaf_memory[9] <= 1;
      stuckIsLeaf_memory[10] <= 1;
      for(stuckIsLeaf_memory_index = 11; stuckIsLeaf_memory_index < 12; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
      stuckIsLeaf_memory[12] <= 1;
      for(stuckIsLeaf_memory_index = 13; stuckIsLeaf_memory_index < 32; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
    end
    else if (processCurrent == 0) begin
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_7_result_0 <= stuckIsLeaf_memory[delete_stuckIsLeaf_7_index_35*1+0];
            stuckIsLeaf_7_finishedAt <= step;
          end
          else if ((stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step)) begin
            stuckIsLeaf_memory[delete_stuckIsLeaf_8_index_36*1+0] <= delete_stuckIsLeaf_8_value_37;
            stuckIsLeaf_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[32*1];
  integer stuckIsFree_11_requestedAt;
  integer stuckIsFree_11_finishedAt;
  integer stuckIsFree_stuckIsFree_11_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  integer stuckIsFree_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_11_finishedAt <= -1;
      stuckIsFree_stuckIsFree_11_returnCode <= 0;
      for(stuckIsFree_memory_index = 0; stuckIsFree_memory_index < 6; stuckIsFree_memory_index = stuckIsFree_memory_index + 1) stuckIsFree_memory[stuckIsFree_memory_index] <= 0;
      stuckIsFree_memory[6] <= 1;
      for(stuckIsFree_memory_index = 7; stuckIsFree_memory_index < 12; stuckIsFree_memory_index = stuckIsFree_memory_index + 1) stuckIsFree_memory[stuckIsFree_memory_index] <= 0;
      stuckIsFree_memory[12] <= 1;
      stuckIsFree_memory[13] <= 1;
      stuckIsFree_memory[14] <= 1;
      stuckIsFree_memory[15] <= 1;
      stuckIsFree_memory[16] <= 1;
      stuckIsFree_memory[17] <= 1;
      stuckIsFree_memory[18] <= 1;
      stuckIsFree_memory[19] <= 1;
      stuckIsFree_memory[20] <= 1;
      stuckIsFree_memory[21] <= 1;
      stuckIsFree_memory[22] <= 1;
      stuckIsFree_memory[23] <= 1;
      stuckIsFree_memory[24] <= 1;
      stuckIsFree_memory[25] <= 1;
      stuckIsFree_memory[26] <= 1;
      stuckIsFree_memory[27] <= 1;
      stuckIsFree_memory[28] <= 1;
      stuckIsFree_memory[29] <= 1;
      stuckIsFree_memory[30] <= 1;
      stuckIsFree_memory[31] <= 1;
    end
    else if (processCurrent == 1) begin
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step)) begin
            stuckIsFree_memory[delete_stuckIsFree_11_index_199*1+0] <= delete_stuckIsFree_11_value_200;
            stuckIsFree_11_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [6-1:0] freeNext_memory[32*1];
  reg [6-1:0] freeNext_freeNext_9_result_0;
  integer freeNext_9_requestedAt;
  integer freeNext_9_finishedAt;
  integer freeNext_freeNext_9_returnCode;
  integer freeNext_10_requestedAt;
  integer freeNext_10_finishedAt;
  integer freeNext_freeNext_10_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  integer freeNext_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_9_result_0 <= 0;
      freeNext_9_finishedAt <= -1;
      freeNext_freeNext_9_returnCode <= 0;
      freeNext_10_finishedAt <= -1;
      freeNext_freeNext_10_returnCode <= 0;
      freeNext_memory[0] <= 6;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 12;
      freeNext_memory[7] <= 8;
      freeNext_memory[8] <= 9;
      freeNext_memory[9] <= 11;
      freeNext_memory[10] <= 9;
      freeNext_memory[11] <= 12;
      freeNext_memory[12] <= 13;
      freeNext_memory[13] <= 14;
      freeNext_memory[14] <= 15;
      freeNext_memory[15] <= 16;
      freeNext_memory[16] <= 17;
      freeNext_memory[17] <= 18;
      freeNext_memory[18] <= 19;
      freeNext_memory[19] <= 20;
      freeNext_memory[20] <= 21;
      freeNext_memory[21] <= 22;
      freeNext_memory[22] <= 23;
      freeNext_memory[23] <= 24;
      freeNext_memory[24] <= 25;
      freeNext_memory[25] <= 26;
      freeNext_memory[26] <= 27;
      freeNext_memory[27] <= 28;
      freeNext_memory[28] <= 29;
      freeNext_memory[29] <= 30;
      freeNext_memory[30] <= 31;
      for(freeNext_memory_index = 31; freeNext_memory_index < 32; freeNext_memory_index = freeNext_memory_index + 1) freeNext_memory[freeNext_memory_index] <= 0;
    end
    else if (processCurrent == 2) begin
      case(freeNext_pc)
        0: begin
          if ((freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step)) begin
            freeNext_freeNext_9_result_0 <= freeNext_memory[delete_freeNext_9_index_196*1+0];
            freeNext_9_finishedAt <= step;
          end
          else if ((freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step)) begin
            freeNext_memory[delete_freeNext_10_index_197*1+0] <= delete_freeNext_10_value_198;
            freeNext_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[32*1];
  reg [3-1:0] stuckSize_stuckSize_5_result_0;
  integer stuckSize_5_requestedAt;
  integer stuckSize_5_finishedAt;
  integer stuckSize_stuckSize_5_returnCode;
  integer stuckSize_6_requestedAt;
  integer stuckSize_6_finishedAt;
  integer stuckSize_stuckSize_6_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  integer stuckSize_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_5_result_0 <= 0;
      stuckSize_5_finishedAt <= -1;
      stuckSize_stuckSize_5_returnCode <= 0;
      stuckSize_6_finishedAt <= -1;
      stuckSize_stuckSize_6_returnCode <= 0;
      stuckSize_memory[0] <= 1;
      stuckSize_memory[1] <= 4;
      stuckSize_memory[2] <= 4;
      stuckSize_memory[3] <= 4;
      stuckSize_memory[4] <= 4;
      stuckSize_memory[5] <= 3;
      stuckSize_memory[6] <= 1;
      stuckSize_memory[7] <= 4;
      stuckSize_memory[8] <= 4;
      stuckSize_memory[9] <= 4;
      stuckSize_memory[10] <= 4;
      stuckSize_memory[11] <= 3;
      stuckSize_memory[12] <= 2;
      for(stuckSize_memory_index = 13; stuckSize_memory_index < 32; stuckSize_memory_index = stuckSize_memory_index + 1) stuckSize_memory[stuckSize_memory_index] <= 0;
    end
    else if (processCurrent == 3) begin
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step)) begin
            stuckSize_stuckSize_5_result_0 <= stuckSize_memory[delete_stuckSize_5_index_32*1+0];
            stuckSize_5_finishedAt <= step;
          end
          else if ((stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step)) begin
            stuckSize_memory[delete_stuckSize_6_index_33*1+0] <= delete_stuckSize_6_value_34;
            stuckSize_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys  process_stuckKeys_0004
  (* ram_style = "block" *)
  reg [8-1:0] stuckKeys_memory[32*4];
  reg [8-1:0] stuckKeys_stuckKeys_1_result_0;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_1;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_2;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_3;
  integer stuckKeys_1_requestedAt;
  integer stuckKeys_1_finishedAt;
  integer stuckKeys_stuckKeys_1_returnCode;
  integer stuckKeys_2_requestedAt;
  integer stuckKeys_2_finishedAt;
  integer stuckKeys_stuckKeys_2_returnCode;
  integer stuckKeys_pc;
  integer stuckKeys_stop;
  integer stuckKeys_returnCode;
  integer stuckKeys_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_pc <= 0;
      stuckKeys_stop <= 0;
      stuckKeys_returnCode <= 0;
      stuckKeys_stuckKeys_1_result_0 <= 0;
      stuckKeys_stuckKeys_1_result_1 <= 0;
      stuckKeys_stuckKeys_1_result_2 <= 0;
      stuckKeys_stuckKeys_1_result_3 <= 0;
      stuckKeys_1_finishedAt <= -1;
      stuckKeys_stuckKeys_1_returnCode <= 0;
      stuckKeys_2_finishedAt <= -1;
      stuckKeys_stuckKeys_2_returnCode <= 0;
      stuckKeys_memory[0] <= 16;
      stuckKeys_memory[1] <= 24;
      stuckKeys_memory[2] <= 24;
      stuckKeys_memory[3] <= 10;
      stuckKeys_memory[4] <= 1;
      stuckKeys_memory[5] <= 2;
      stuckKeys_memory[6] <= 3;
      stuckKeys_memory[7] <= 4;
      stuckKeys_memory[8] <= 29;
      stuckKeys_memory[9] <= 30;
      stuckKeys_memory[10] <= 31;
      stuckKeys_memory[11] <= 32;
      stuckKeys_memory[12] <= 5;
      stuckKeys_memory[13] <= 6;
      stuckKeys_memory[14] <= 7;
      stuckKeys_memory[15] <= 8;
      stuckKeys_memory[16] <= 9;
      stuckKeys_memory[17] <= 10;
      stuckKeys_memory[18] <= 11;
      stuckKeys_memory[19] <= 12;
      stuckKeys_memory[20] <= 4;
      stuckKeys_memory[21] <= 8;
      stuckKeys_memory[22] <= 12;
      for(stuckKeys_memory_index = 23; stuckKeys_memory_index < 24; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
      stuckKeys_memory[24] <= 28;
      stuckKeys_memory[25] <= 28;
      stuckKeys_memory[26] <= 26;
      stuckKeys_memory[27] <= 26;
      stuckKeys_memory[28] <= 13;
      stuckKeys_memory[29] <= 14;
      stuckKeys_memory[30] <= 15;
      stuckKeys_memory[31] <= 16;
      stuckKeys_memory[32] <= 17;
      stuckKeys_memory[33] <= 18;
      stuckKeys_memory[34] <= 19;
      stuckKeys_memory[35] <= 20;
      stuckKeys_memory[36] <= 25;
      stuckKeys_memory[37] <= 26;
      stuckKeys_memory[38] <= 27;
      stuckKeys_memory[39] <= 28;
      stuckKeys_memory[40] <= 21;
      stuckKeys_memory[41] <= 22;
      stuckKeys_memory[42] <= 23;
      stuckKeys_memory[43] <= 24;
      stuckKeys_memory[44] <= 20;
      stuckKeys_memory[45] <= 24;
      stuckKeys_memory[46] <= 28;
      for(stuckKeys_memory_index = 47; stuckKeys_memory_index < 48; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
      stuckKeys_memory[48] <= 27;
      stuckKeys_memory[49] <= 28;
      for(stuckKeys_memory_index = 50; stuckKeys_memory_index < 128; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
    end
    else if (processCurrent == 4) begin
      case(stuckKeys_pc)
        0: begin
          if ((stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step)) begin
            stuckKeys_stuckKeys_1_result_0 <= stuckKeys_memory[delete_stuckKeys_1_index_20*4+0];
            stuckKeys_stuckKeys_1_result_1 <= stuckKeys_memory[delete_stuckKeys_1_index_20*4+1];
            stuckKeys_stuckKeys_1_result_2 <= stuckKeys_memory[delete_stuckKeys_1_index_20*4+2];
            stuckKeys_stuckKeys_1_result_3 <= stuckKeys_memory[delete_stuckKeys_1_index_20*4+3];
            stuckKeys_1_finishedAt <= step;
          end
          else if ((stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step)) begin
            stuckKeys_memory[delete_stuckKeys_2_index_21*4+0] <= delete_stuckKeys_2_value_22;
            stuckKeys_memory[delete_stuckKeys_2_index_21*4+1] <= delete_stuckKeys_2_value_23;
            stuckKeys_memory[delete_stuckKeys_2_index_21*4+2] <= delete_stuckKeys_2_value_24;
            stuckKeys_memory[delete_stuckKeys_2_index_21*4+3] <= delete_stuckKeys_2_value_25;
            stuckKeys_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_stop <= 1;
      endcase
    end
  end
  // Process: stuckData  process_stuckData_0005
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_memory[32*4];
  reg [8-1:0] stuckData_stuckData_3_result_0;
  reg [8-1:0] stuckData_stuckData_3_result_1;
  reg [8-1:0] stuckData_stuckData_3_result_2;
  reg [8-1:0] stuckData_stuckData_3_result_3;
  integer stuckData_3_requestedAt;
  integer stuckData_3_finishedAt;
  integer stuckData_stuckData_3_returnCode;
  integer stuckData_4_requestedAt;
  integer stuckData_4_finishedAt;
  integer stuckData_stuckData_4_returnCode;
  integer stuckData_pc;
  integer stuckData_stop;
  integer stuckData_returnCode;
  integer stuckData_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_pc <= 0;
      stuckData_stop <= 0;
      stuckData_returnCode <= 0;
      stuckData_stuckData_3_result_0 <= 0;
      stuckData_stuckData_3_result_1 <= 0;
      stuckData_stuckData_3_result_2 <= 0;
      stuckData_stuckData_3_result_3 <= 0;
      stuckData_3_finishedAt <= -1;
      stuckData_stuckData_3_returnCode <= 0;
      stuckData_4_finishedAt <= -1;
      stuckData_stuckData_4_returnCode <= 0;
      stuckData_memory[0] <= 5;
      stuckData_memory[1] <= 11;
      stuckData_memory[2] <= 6;
      stuckData_memory[3] <= 2;
      stuckData_memory[4] <= 2;
      stuckData_memory[5] <= 3;
      stuckData_memory[6] <= 4;
      stuckData_memory[7] <= 5;
      stuckData_memory[8] <= 30;
      stuckData_memory[9] <= 31;
      stuckData_memory[10] <= 32;
      stuckData_memory[11] <= 33;
      stuckData_memory[12] <= 6;
      stuckData_memory[13] <= 7;
      stuckData_memory[14] <= 8;
      stuckData_memory[15] <= 9;
      stuckData_memory[16] <= 10;
      stuckData_memory[17] <= 11;
      stuckData_memory[18] <= 12;
      stuckData_memory[19] <= 13;
      stuckData_memory[20] <= 1;
      stuckData_memory[21] <= 3;
      stuckData_memory[22] <= 4;
      stuckData_memory[23] <= 7;
      stuckData_memory[24] <= 9;
      stuckData_memory[25] <= 2;
      stuckData_memory[26] <= 2;
      stuckData_memory[27] <= 2;
      stuckData_memory[28] <= 14;
      stuckData_memory[29] <= 15;
      stuckData_memory[30] <= 16;
      stuckData_memory[31] <= 17;
      stuckData_memory[32] <= 18;
      stuckData_memory[33] <= 19;
      stuckData_memory[34] <= 20;
      stuckData_memory[35] <= 21;
      stuckData_memory[36] <= 26;
      stuckData_memory[37] <= 27;
      stuckData_memory[38] <= 28;
      stuckData_memory[39] <= 29;
      stuckData_memory[40] <= 22;
      stuckData_memory[41] <= 23;
      stuckData_memory[42] <= 24;
      stuckData_memory[43] <= 25;
      stuckData_memory[44] <= 8;
      stuckData_memory[45] <= 10;
      stuckData_memory[46] <= 9;
      stuckData_memory[47] <= 2;
      stuckData_memory[48] <= 28;
      stuckData_memory[49] <= 29;
      for(stuckData_memory_index = 50; stuckData_memory_index < 128; stuckData_memory_index = stuckData_memory_index + 1) stuckData_memory[stuckData_memory_index] <= 0;
    end
    else if (processCurrent == 5) begin
      case(stuckData_pc)
        0: begin
          if ((stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step)) begin
            stuckData_stuckData_3_result_0 <= stuckData_memory[delete_stuckData_3_index_26*4+0];
            stuckData_stuckData_3_result_1 <= stuckData_memory[delete_stuckData_3_index_26*4+1];
            stuckData_stuckData_3_result_2 <= stuckData_memory[delete_stuckData_3_index_26*4+2];
            stuckData_stuckData_3_result_3 <= stuckData_memory[delete_stuckData_3_index_26*4+3];
            stuckData_3_finishedAt <= step;
          end
          else if ((stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step)) begin
            stuckData_memory[delete_stuckData_4_index_27*4+0] <= delete_stuckData_4_value_28;
            stuckData_memory[delete_stuckData_4_index_27*4+1] <= delete_stuckData_4_value_29;
            stuckData_memory[delete_stuckData_4_index_27*4+2] <= delete_stuckData_4_value_30;
            stuckData_memory[delete_stuckData_4_index_27*4+3] <= delete_stuckData_4_value_31;
            stuckData_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_stop <= 1;
      endcase
    end
  end
  // Process: delete  process_delete_0006
  reg [6-1:0] delete_index_0;
  reg [3-1:0] delete_size_1;
  reg [1-1:0] delete_isLeaf_2;
  reg [6-1:0] delete_nextFree_3;
  reg [8-1:0] delete_Key_0_4;
  reg [1-1:0] delete_KeyCompares_0_5;
  reg [3-1:0] delete_KeyCollapse_0_6;
  reg [8-1:0] delete_Data_0_7;
  reg [8-1:0] delete_Key_1_8;
  reg [1-1:0] delete_KeyCompares_1_9;
  reg [3-1:0] delete_KeyCollapse_1_10;
  reg [8-1:0] delete_Data_1_11;
  reg [8-1:0] delete_Key_2_12;
  reg [1-1:0] delete_KeyCompares_2_13;
  reg [3-1:0] delete_KeyCollapse_2_14;
  reg [8-1:0] delete_Data_2_15;
  reg [8-1:0] delete_Key_3_16;
  reg [1-1:0] delete_KeyCompares_3_17;
  reg [3-1:0] delete_KeyCollapse_3_18;
  reg [8-1:0] delete_Data_3_19;
  reg [5-1:0] delete_stuckKeys_1_index_20;
  reg [5-1:0] delete_stuckKeys_2_index_21;
  reg [8-1:0] delete_stuckKeys_2_value_22;
  reg [8-1:0] delete_stuckKeys_2_value_23;
  reg [8-1:0] delete_stuckKeys_2_value_24;
  reg [8-1:0] delete_stuckKeys_2_value_25;
  reg [5-1:0] delete_stuckData_3_index_26;
  reg [5-1:0] delete_stuckData_4_index_27;
  reg [8-1:0] delete_stuckData_4_value_28;
  reg [8-1:0] delete_stuckData_4_value_29;
  reg [8-1:0] delete_stuckData_4_value_30;
  reg [8-1:0] delete_stuckData_4_value_31;
  reg [5-1:0] delete_stuckSize_5_index_32;
  reg [5-1:0] delete_stuckSize_6_index_33;
  reg [3-1:0] delete_stuckSize_6_value_34;
  reg [5-1:0] delete_stuckIsLeaf_7_index_35;
  reg [5-1:0] delete_stuckIsLeaf_8_index_36;
  reg [1-1:0] delete_stuckIsLeaf_8_value_37;
  reg [1-1:0] delete_Found_38;
  reg [8-1:0] delete_Key_39;
  reg [8-1:0] delete_FoundKey_40;
  reg [8-1:0] delete_Data_41;
  reg [6-1:0] delete_BtreeIndex_42;
  reg [3-1:0] delete_StuckIndex_43;
  reg [1-1:0] delete_MergeSuccess_44;
  reg [6-1:0] delete_i_45;
  reg [8-1:0] delete_k_46;
  reg [1-1:0] delete_l_47;
  reg [6-1:0] delete_index_48;
  reg [3-1:0] delete_size_49;
  reg [1-1:0] delete_isLeaf_50;
  reg [6-1:0] delete_nextFree_51;
  reg [8-1:0] delete_Key_0_52;
  reg [1-1:0] delete_KeyCompares_0_53;
  reg [3-1:0] delete_KeyCollapse_0_54;
  reg [8-1:0] delete_Data_0_55;
  reg [8-1:0] delete_Key_1_56;
  reg [1-1:0] delete_KeyCompares_1_57;
  reg [3-1:0] delete_KeyCollapse_1_58;
  reg [8-1:0] delete_Data_1_59;
  reg [8-1:0] delete_Key_2_60;
  reg [1-1:0] delete_KeyCompares_2_61;
  reg [3-1:0] delete_KeyCollapse_2_62;
  reg [8-1:0] delete_Data_2_63;
  reg [8-1:0] delete_Key_3_64;
  reg [1-1:0] delete_KeyCompares_3_65;
  reg [3-1:0] delete_KeyCollapse_3_66;
  reg [8-1:0] delete_Data_3_67;
  reg [1-1:0] delete_Found_68;
  reg [8-1:0] delete_Key_69;
  reg [8-1:0] delete_FoundKey_70;
  reg [8-1:0] delete_Data_71;
  reg [6-1:0] delete_BtreeIndex_72;
  reg [3-1:0] delete_StuckIndex_73;
  reg [1-1:0] delete_MergeSuccess_74;
  reg [6-1:0] delete_index_75;
  reg [3-1:0] delete_size_76;
  reg [1-1:0] delete_isLeaf_77;
  reg [6-1:0] delete_nextFree_78;
  reg [8-1:0] delete_Key_0_79;
  reg [1-1:0] delete_KeyCompares_0_80;
  reg [3-1:0] delete_KeyCollapse_0_81;
  reg [8-1:0] delete_Data_0_82;
  reg [8-1:0] delete_Key_1_83;
  reg [1-1:0] delete_KeyCompares_1_84;
  reg [3-1:0] delete_KeyCollapse_1_85;
  reg [8-1:0] delete_Data_1_86;
  reg [8-1:0] delete_Key_2_87;
  reg [1-1:0] delete_KeyCompares_2_88;
  reg [3-1:0] delete_KeyCollapse_2_89;
  reg [8-1:0] delete_Data_2_90;
  reg [8-1:0] delete_Key_3_91;
  reg [1-1:0] delete_KeyCompares_3_92;
  reg [3-1:0] delete_KeyCollapse_3_93;
  reg [8-1:0] delete_Data_3_94;
  reg [1-1:0] delete_Found_95;
  reg [8-1:0] delete_Key_96;
  reg [8-1:0] delete_FoundKey_97;
  reg [8-1:0] delete_Data_98;
  reg [6-1:0] delete_BtreeIndex_99;
  reg [3-1:0] delete_StuckIndex_100;
  reg [1-1:0] delete_MergeSuccess_101;
  reg [6-1:0] delete_position_102;
  reg [3-1:0] delete_index_103;
  reg [3-1:0] delete_index1_104;
  reg [1-1:0] delete_within_105;
  reg [1-1:0] delete_isLeaf_106;
  reg [6-1:0] delete_index_107;
  reg [3-1:0] delete_size_108;
  reg [1-1:0] delete_isLeaf_109;
  reg [6-1:0] delete_nextFree_110;
  reg [8-1:0] delete_Key_0_111;
  reg [1-1:0] delete_KeyCompares_0_112;
  reg [3-1:0] delete_KeyCollapse_0_113;
  reg [8-1:0] delete_Data_0_114;
  reg [8-1:0] delete_Key_1_115;
  reg [1-1:0] delete_KeyCompares_1_116;
  reg [3-1:0] delete_KeyCollapse_1_117;
  reg [8-1:0] delete_Data_1_118;
  reg [8-1:0] delete_Key_2_119;
  reg [1-1:0] delete_KeyCompares_2_120;
  reg [3-1:0] delete_KeyCollapse_2_121;
  reg [8-1:0] delete_Data_2_122;
  reg [8-1:0] delete_Key_3_123;
  reg [1-1:0] delete_KeyCompares_3_124;
  reg [3-1:0] delete_KeyCollapse_3_125;
  reg [8-1:0] delete_Data_3_126;
  reg [1-1:0] delete_Found_127;
  reg [8-1:0] delete_Key_128;
  reg [8-1:0] delete_FoundKey_129;
  reg [8-1:0] delete_Data_130;
  reg [6-1:0] delete_BtreeIndex_131;
  reg [3-1:0] delete_StuckIndex_132;
  reg [1-1:0] delete_MergeSuccess_133;
  reg [6-1:0] delete_index_134;
  reg [3-1:0] delete_size_135;
  reg [1-1:0] delete_isLeaf_136;
  reg [6-1:0] delete_nextFree_137;
  reg [8-1:0] delete_Key_0_138;
  reg [1-1:0] delete_KeyCompares_0_139;
  reg [3-1:0] delete_KeyCollapse_0_140;
  reg [8-1:0] delete_Data_0_141;
  reg [8-1:0] delete_Key_1_142;
  reg [1-1:0] delete_KeyCompares_1_143;
  reg [3-1:0] delete_KeyCollapse_1_144;
  reg [8-1:0] delete_Data_1_145;
  reg [8-1:0] delete_Key_2_146;
  reg [1-1:0] delete_KeyCompares_2_147;
  reg [3-1:0] delete_KeyCollapse_2_148;
  reg [8-1:0] delete_Data_2_149;
  reg [8-1:0] delete_Key_3_150;
  reg [1-1:0] delete_KeyCompares_3_151;
  reg [3-1:0] delete_KeyCollapse_3_152;
  reg [8-1:0] delete_Data_3_153;
  reg [1-1:0] delete_Found_154;
  reg [8-1:0] delete_Key_155;
  reg [8-1:0] delete_FoundKey_156;
  reg [8-1:0] delete_Data_157;
  reg [6-1:0] delete_BtreeIndex_158;
  reg [3-1:0] delete_StuckIndex_159;
  reg [1-1:0] delete_MergeSuccess_160;
  reg [6-1:0] delete_index_161;
  reg [3-1:0] delete_size_162;
  reg [1-1:0] delete_isLeaf_163;
  reg [6-1:0] delete_nextFree_164;
  reg [8-1:0] delete_Key_0_165;
  reg [1-1:0] delete_KeyCompares_0_166;
  reg [3-1:0] delete_KeyCollapse_0_167;
  reg [8-1:0] delete_Data_0_168;
  reg [8-1:0] delete_Key_1_169;
  reg [1-1:0] delete_KeyCompares_1_170;
  reg [3-1:0] delete_KeyCollapse_1_171;
  reg [8-1:0] delete_Data_1_172;
  reg [8-1:0] delete_Key_2_173;
  reg [1-1:0] delete_KeyCompares_2_174;
  reg [3-1:0] delete_KeyCollapse_2_175;
  reg [8-1:0] delete_Data_2_176;
  reg [8-1:0] delete_Key_3_177;
  reg [1-1:0] delete_KeyCompares_3_178;
  reg [3-1:0] delete_KeyCollapse_3_179;
  reg [8-1:0] delete_Data_3_180;
  reg [1-1:0] delete_Found_181;
  reg [8-1:0] delete_Key_182;
  reg [8-1:0] delete_FoundKey_183;
  reg [8-1:0] delete_Data_184;
  reg [6-1:0] delete_BtreeIndex_185;
  reg [3-1:0] delete_StuckIndex_186;
  reg [1-1:0] delete_MergeSuccess_187;
  reg [8-1:0] delete_childKey_188;
  reg [6-1:0] delete_childData_189;
  reg [6-1:0] delete_indexLeft_190;
  reg [6-1:0] delete_indexRight_191;
  reg [8-1:0] delete_midKey_192;
  reg [1-1:0] delete_success_193;
  reg [1-1:0] delete_test_194;
  reg [6-1:0] delete_next_195;
  reg [5-1:0] delete_freeNext_9_index_196;
  reg [5-1:0] delete_freeNext_10_index_197;
  reg [6-1:0] delete_freeNext_10_value_198;
  reg [5-1:0] delete_stuckIsFree_11_index_199;
  reg [1-1:0] delete_stuckIsFree_11_value_200;
  reg [6-1:0] delete_root_201;
  reg [1-1:0] delete_isFree_202;
  reg [6-1:0] delete_next_203;
  reg [6-1:0] delete_root_204;
  reg [1-1:0] delete_isFree_205;
  reg [6-1:0] delete_index_206;
  reg [3-1:0] delete_size_207;
  reg [1-1:0] delete_isLeaf_208;
  reg [6-1:0] delete_nextFree_209;
  reg [8-1:0] delete_Key_0_210;
  reg [1-1:0] delete_KeyCompares_0_211;
  reg [3-1:0] delete_KeyCollapse_0_212;
  reg [8-1:0] delete_Data_0_213;
  reg [8-1:0] delete_Key_1_214;
  reg [1-1:0] delete_KeyCompares_1_215;
  reg [3-1:0] delete_KeyCollapse_1_216;
  reg [8-1:0] delete_Data_1_217;
  reg [8-1:0] delete_Key_2_218;
  reg [1-1:0] delete_KeyCompares_2_219;
  reg [3-1:0] delete_KeyCollapse_2_220;
  reg [8-1:0] delete_Data_2_221;
  reg [8-1:0] delete_Key_3_222;
  reg [1-1:0] delete_KeyCompares_3_223;
  reg [3-1:0] delete_KeyCollapse_3_224;
  reg [8-1:0] delete_Data_3_225;
  reg [1-1:0] delete_Found_226;
  reg [8-1:0] delete_Key_227;
  reg [8-1:0] delete_FoundKey_228;
  reg [8-1:0] delete_Data_229;
  reg [6-1:0] delete_BtreeIndex_230;
  reg [3-1:0] delete_StuckIndex_231;
  reg [1-1:0] delete_MergeSuccess_232;
  reg [6-1:0] delete_index_233;
  reg [3-1:0] delete_size_234;
  reg [1-1:0] delete_isLeaf_235;
  reg [6-1:0] delete_nextFree_236;
  reg [8-1:0] delete_Key_0_237;
  reg [1-1:0] delete_KeyCompares_0_238;
  reg [3-1:0] delete_KeyCollapse_0_239;
  reg [8-1:0] delete_Data_0_240;
  reg [8-1:0] delete_Key_1_241;
  reg [1-1:0] delete_KeyCompares_1_242;
  reg [3-1:0] delete_KeyCollapse_1_243;
  reg [8-1:0] delete_Data_1_244;
  reg [8-1:0] delete_Key_2_245;
  reg [1-1:0] delete_KeyCompares_2_246;
  reg [3-1:0] delete_KeyCollapse_2_247;
  reg [8-1:0] delete_Data_2_248;
  reg [8-1:0] delete_Key_3_249;
  reg [1-1:0] delete_KeyCompares_3_250;
  reg [3-1:0] delete_KeyCollapse_3_251;
  reg [8-1:0] delete_Data_3_252;
  reg [1-1:0] delete_Found_253;
  reg [8-1:0] delete_Key_254;
  reg [8-1:0] delete_FoundKey_255;
  reg [8-1:0] delete_Data_256;
  reg [6-1:0] delete_BtreeIndex_257;
  reg [3-1:0] delete_StuckIndex_258;
  reg [1-1:0] delete_MergeSuccess_259;
  reg [6-1:0] delete_index_260;
  reg [3-1:0] delete_size_261;
  reg [1-1:0] delete_isLeaf_262;
  reg [6-1:0] delete_nextFree_263;
  reg [8-1:0] delete_Key_0_264;
  reg [1-1:0] delete_KeyCompares_0_265;
  reg [3-1:0] delete_KeyCollapse_0_266;
  reg [8-1:0] delete_Data_0_267;
  reg [8-1:0] delete_Key_1_268;
  reg [1-1:0] delete_KeyCompares_1_269;
  reg [3-1:0] delete_KeyCollapse_1_270;
  reg [8-1:0] delete_Data_1_271;
  reg [8-1:0] delete_Key_2_272;
  reg [1-1:0] delete_KeyCompares_2_273;
  reg [3-1:0] delete_KeyCollapse_2_274;
  reg [8-1:0] delete_Data_2_275;
  reg [8-1:0] delete_Key_3_276;
  reg [1-1:0] delete_KeyCompares_3_277;
  reg [3-1:0] delete_KeyCollapse_3_278;
  reg [8-1:0] delete_Data_3_279;
  reg [1-1:0] delete_Found_280;
  reg [8-1:0] delete_Key_281;
  reg [8-1:0] delete_FoundKey_282;
  reg [8-1:0] delete_Data_283;
  reg [6-1:0] delete_BtreeIndex_284;
  reg [3-1:0] delete_StuckIndex_285;
  reg [1-1:0] delete_MergeSuccess_286;
  reg [8-1:0] delete_childKey_287;
  reg [3-1:0] delete_leftChild_288;
  reg [3-1:0] delete_rightChild_289;
  reg [6-1:0] delete_childData_290;
  reg [6-1:0] delete_indexLeft_291;
  reg [6-1:0] delete_indexRight_292;
  reg [8-1:0] delete_midKey_293;
  reg [1-1:0] delete_success_294;
  reg [1-1:0] delete_test_295;
  reg [6-1:0] delete_next_296;
  reg [6-1:0] delete_root_297;
  reg [1-1:0] delete_isFree_298;
  reg [6-1:0] delete_next_299;
  reg [6-1:0] delete_root_300;
  reg [1-1:0] delete_isFree_301;
  reg [6-1:0] delete_index_302;
  reg [3-1:0] delete_size_303;
  reg [1-1:0] delete_isLeaf_304;
  reg [6-1:0] delete_nextFree_305;
  reg [8-1:0] delete_Key_0_306;
  reg [1-1:0] delete_KeyCompares_0_307;
  reg [3-1:0] delete_KeyCollapse_0_308;
  reg [8-1:0] delete_Data_0_309;
  reg [8-1:0] delete_Key_1_310;
  reg [1-1:0] delete_KeyCompares_1_311;
  reg [3-1:0] delete_KeyCollapse_1_312;
  reg [8-1:0] delete_Data_1_313;
  reg [8-1:0] delete_Key_2_314;
  reg [1-1:0] delete_KeyCompares_2_315;
  reg [3-1:0] delete_KeyCollapse_2_316;
  reg [8-1:0] delete_Data_2_317;
  reg [8-1:0] delete_Key_3_318;
  reg [1-1:0] delete_KeyCompares_3_319;
  reg [3-1:0] delete_KeyCollapse_3_320;
  reg [8-1:0] delete_Data_3_321;
  reg [1-1:0] delete_Found_322;
  reg [8-1:0] delete_Key_323;
  reg [8-1:0] delete_FoundKey_324;
  reg [8-1:0] delete_Data_325;
  reg [6-1:0] delete_BtreeIndex_326;
  reg [3-1:0] delete_StuckIndex_327;
  reg [1-1:0] delete_MergeSuccess_328;
  reg [6-1:0] delete_index_329;
  reg [3-1:0] delete_size_330;
  reg [1-1:0] delete_isLeaf_331;
  reg [6-1:0] delete_nextFree_332;
  reg [8-1:0] delete_Key_0_333;
  reg [1-1:0] delete_KeyCompares_0_334;
  reg [3-1:0] delete_KeyCollapse_0_335;
  reg [8-1:0] delete_Data_0_336;
  reg [8-1:0] delete_Key_1_337;
  reg [1-1:0] delete_KeyCompares_1_338;
  reg [3-1:0] delete_KeyCollapse_1_339;
  reg [8-1:0] delete_Data_1_340;
  reg [8-1:0] delete_Key_2_341;
  reg [1-1:0] delete_KeyCompares_2_342;
  reg [3-1:0] delete_KeyCollapse_2_343;
  reg [8-1:0] delete_Data_2_344;
  reg [8-1:0] delete_Key_3_345;
  reg [1-1:0] delete_KeyCompares_3_346;
  reg [3-1:0] delete_KeyCollapse_3_347;
  reg [8-1:0] delete_Data_3_348;
  reg [1-1:0] delete_Found_349;
  reg [8-1:0] delete_Key_350;
  reg [8-1:0] delete_FoundKey_351;
  reg [8-1:0] delete_Data_352;
  reg [6-1:0] delete_BtreeIndex_353;
  reg [3-1:0] delete_StuckIndex_354;
  reg [1-1:0] delete_MergeSuccess_355;
  reg [8-1:0] delete_childKey_356;
  reg [3-1:0] delete_size_357;
  reg [6-1:0] delete_childData_358;
  reg [6-1:0] delete_indexLeft_359;
  reg [6-1:0] delete_indexRight_360;
  reg [8-1:0] delete_midKey_361;
  reg [1-1:0] delete_success_362;
  reg [1-1:0] delete_test_363;
  reg [6-1:0] delete_next_364;
  reg [6-1:0] delete_root_365;
  reg [1-1:0] delete_isFree_366;
  reg [6-1:0] delete_index_367;
  reg [3-1:0] delete_size_368;
  reg [1-1:0] delete_isLeaf_369;
  reg [6-1:0] delete_nextFree_370;
  reg [8-1:0] delete_Key_0_371;
  reg [1-1:0] delete_KeyCompares_0_372;
  reg [3-1:0] delete_KeyCollapse_0_373;
  reg [8-1:0] delete_Data_0_374;
  reg [8-1:0] delete_Key_1_375;
  reg [1-1:0] delete_KeyCompares_1_376;
  reg [3-1:0] delete_KeyCollapse_1_377;
  reg [8-1:0] delete_Data_1_378;
  reg [8-1:0] delete_Key_2_379;
  reg [1-1:0] delete_KeyCompares_2_380;
  reg [3-1:0] delete_KeyCollapse_2_381;
  reg [8-1:0] delete_Data_2_382;
  reg [8-1:0] delete_Key_3_383;
  reg [1-1:0] delete_KeyCompares_3_384;
  reg [3-1:0] delete_KeyCollapse_3_385;
  reg [8-1:0] delete_Data_3_386;
  reg [1-1:0] delete_Found_387;
  reg [8-1:0] delete_Key_388;
  reg [8-1:0] delete_FoundKey_389;
  reg [8-1:0] delete_Data_390;
  reg [6-1:0] delete_BtreeIndex_391;
  reg [3-1:0] delete_StuckIndex_392;
  reg [1-1:0] delete_MergeSuccess_393;
  reg [6-1:0] delete_index_394;
  reg [3-1:0] delete_size_395;
  reg [1-1:0] delete_isLeaf_396;
  reg [6-1:0] delete_nextFree_397;
  reg [8-1:0] delete_Key_0_398;
  reg [1-1:0] delete_KeyCompares_0_399;
  reg [3-1:0] delete_KeyCollapse_0_400;
  reg [8-1:0] delete_Data_0_401;
  reg [8-1:0] delete_Key_1_402;
  reg [1-1:0] delete_KeyCompares_1_403;
  reg [3-1:0] delete_KeyCollapse_1_404;
  reg [8-1:0] delete_Data_1_405;
  reg [8-1:0] delete_Key_2_406;
  reg [1-1:0] delete_KeyCompares_2_407;
  reg [3-1:0] delete_KeyCollapse_2_408;
  reg [8-1:0] delete_Data_2_409;
  reg [8-1:0] delete_Key_3_410;
  reg [1-1:0] delete_KeyCompares_3_411;
  reg [3-1:0] delete_KeyCollapse_3_412;
  reg [8-1:0] delete_Data_3_413;
  reg [1-1:0] delete_Found_414;
  reg [8-1:0] delete_Key_415;
  reg [8-1:0] delete_FoundKey_416;
  reg [8-1:0] delete_Data_417;
  reg [6-1:0] delete_BtreeIndex_418;
  reg [3-1:0] delete_StuckIndex_419;
  reg [1-1:0] delete_MergeSuccess_420;
  reg [8-1:0] delete_childKey_421;
  reg [3-1:0] delete_size_422;
  reg [6-1:0] delete_childData_423;
  reg [6-1:0] delete_indexLeft_424;
  reg [6-1:0] delete_indexRight_425;
  reg [8-1:0] delete_midKey_426;
  reg [1-1:0] delete_success_427;
  reg [1-1:0] delete_test_428;
  reg [6-1:0] delete_next_429;
  reg [6-1:0] delete_root_430;
  reg [1-1:0] delete_isFree_431;
  reg [6-1:0] delete_index_432;
  reg [3-1:0] delete_size_433;
  reg [1-1:0] delete_isLeaf_434;
  reg [6-1:0] delete_nextFree_435;
  reg [8-1:0] delete_Key_0_436;
  reg [1-1:0] delete_KeyCompares_0_437;
  reg [3-1:0] delete_KeyCollapse_0_438;
  reg [8-1:0] delete_Data_0_439;
  reg [8-1:0] delete_Key_1_440;
  reg [1-1:0] delete_KeyCompares_1_441;
  reg [3-1:0] delete_KeyCollapse_1_442;
  reg [8-1:0] delete_Data_1_443;
  reg [8-1:0] delete_Key_2_444;
  reg [1-1:0] delete_KeyCompares_2_445;
  reg [3-1:0] delete_KeyCollapse_2_446;
  reg [8-1:0] delete_Data_2_447;
  reg [8-1:0] delete_Key_3_448;
  reg [1-1:0] delete_KeyCompares_3_449;
  reg [3-1:0] delete_KeyCollapse_3_450;
  reg [8-1:0] delete_Data_3_451;
  reg [1-1:0] delete_Found_452;
  reg [8-1:0] delete_Key_453;
  reg [8-1:0] delete_FoundKey_454;
  reg [8-1:0] delete_Data_455;
  reg [6-1:0] delete_BtreeIndex_456;
  reg [3-1:0] delete_StuckIndex_457;
  reg [1-1:0] delete_MergeSuccess_458;
  reg [6-1:0] delete_index_459;
  reg [3-1:0] delete_size_460;
  reg [1-1:0] delete_isLeaf_461;
  reg [6-1:0] delete_nextFree_462;
  reg [8-1:0] delete_Key_0_463;
  reg [1-1:0] delete_KeyCompares_0_464;
  reg [3-1:0] delete_KeyCollapse_0_465;
  reg [8-1:0] delete_Data_0_466;
  reg [8-1:0] delete_Key_1_467;
  reg [1-1:0] delete_KeyCompares_1_468;
  reg [3-1:0] delete_KeyCollapse_1_469;
  reg [8-1:0] delete_Data_1_470;
  reg [8-1:0] delete_Key_2_471;
  reg [1-1:0] delete_KeyCompares_2_472;
  reg [3-1:0] delete_KeyCollapse_2_473;
  reg [8-1:0] delete_Data_2_474;
  reg [8-1:0] delete_Key_3_475;
  reg [1-1:0] delete_KeyCompares_3_476;
  reg [3-1:0] delete_KeyCollapse_3_477;
  reg [8-1:0] delete_Data_3_478;
  reg [1-1:0] delete_Found_479;
  reg [8-1:0] delete_Key_480;
  reg [8-1:0] delete_FoundKey_481;
  reg [8-1:0] delete_Data_482;
  reg [6-1:0] delete_BtreeIndex_483;
  reg [3-1:0] delete_StuckIndex_484;
  reg [1-1:0] delete_MergeSuccess_485;
  reg [8-1:0] delete_childKey_486;
  reg [6-1:0] delete_childData_487;
  reg [6-1:0] delete_indexLeft_488;
  reg [6-1:0] delete_indexRight_489;
  reg [8-1:0] delete_midKey_490;
  reg [1-1:0] delete_success_491;
  reg [1-1:0] delete_test_492;
  reg [6-1:0] delete_next_493;
  reg [6-1:0] delete_root_494;
  reg [1-1:0] delete_isFree_495;
  reg [6-1:0] delete_index_496;
  reg [3-1:0] delete_size_497;
  reg [1-1:0] delete_isLeaf_498;
  reg [6-1:0] delete_nextFree_499;
  reg [8-1:0] delete_Key_0_500;
  reg [1-1:0] delete_KeyCompares_0_501;
  reg [3-1:0] delete_KeyCollapse_0_502;
  reg [8-1:0] delete_Data_0_503;
  reg [8-1:0] delete_Key_1_504;
  reg [1-1:0] delete_KeyCompares_1_505;
  reg [3-1:0] delete_KeyCollapse_1_506;
  reg [8-1:0] delete_Data_1_507;
  reg [8-1:0] delete_Key_2_508;
  reg [1-1:0] delete_KeyCompares_2_509;
  reg [3-1:0] delete_KeyCollapse_2_510;
  reg [8-1:0] delete_Data_2_511;
  reg [8-1:0] delete_Key_3_512;
  reg [1-1:0] delete_KeyCompares_3_513;
  reg [3-1:0] delete_KeyCollapse_3_514;
  reg [8-1:0] delete_Data_3_515;
  reg [1-1:0] delete_Found_516;
  reg [8-1:0] delete_Key_517;
  reg [8-1:0] delete_FoundKey_518;
  reg [8-1:0] delete_Data_519;
  reg [6-1:0] delete_BtreeIndex_520;
  reg [3-1:0] delete_StuckIndex_521;
  reg [1-1:0] delete_MergeSuccess_522;
  reg [6-1:0] delete_index_523;
  reg [3-1:0] delete_size_524;
  reg [1-1:0] delete_isLeaf_525;
  reg [6-1:0] delete_nextFree_526;
  reg [8-1:0] delete_Key_0_527;
  reg [1-1:0] delete_KeyCompares_0_528;
  reg [3-1:0] delete_KeyCollapse_0_529;
  reg [8-1:0] delete_Data_0_530;
  reg [8-1:0] delete_Key_1_531;
  reg [1-1:0] delete_KeyCompares_1_532;
  reg [3-1:0] delete_KeyCollapse_1_533;
  reg [8-1:0] delete_Data_1_534;
  reg [8-1:0] delete_Key_2_535;
  reg [1-1:0] delete_KeyCompares_2_536;
  reg [3-1:0] delete_KeyCollapse_2_537;
  reg [8-1:0] delete_Data_2_538;
  reg [8-1:0] delete_Key_3_539;
  reg [1-1:0] delete_KeyCompares_3_540;
  reg [3-1:0] delete_KeyCollapse_3_541;
  reg [8-1:0] delete_Data_3_542;
  reg [1-1:0] delete_Found_543;
  reg [8-1:0] delete_Key_544;
  reg [8-1:0] delete_FoundKey_545;
  reg [8-1:0] delete_Data_546;
  reg [6-1:0] delete_BtreeIndex_547;
  reg [3-1:0] delete_StuckIndex_548;
  reg [1-1:0] delete_MergeSuccess_549;
  reg [8-1:0] delete_childKey_550;
  reg [3-1:0] delete_leftChild_551;
  reg [3-1:0] delete_rightChild_552;
  reg [6-1:0] delete_childData_553;
  reg [6-1:0] delete_indexLeft_554;
  reg [6-1:0] delete_indexRight_555;
  reg [8-1:0] delete_midKey_556;
  reg [1-1:0] delete_success_557;
  reg [1-1:0] delete_test_558;
  reg [6-1:0] delete_next_559;
  reg [6-1:0] delete_root_560;
  reg [1-1:0] delete_isFree_561;
  reg [6-1:0] delete_index_562;
  reg [3-1:0] delete_size_563;
  reg [1-1:0] delete_isLeaf_564;
  reg [6-1:0] delete_nextFree_565;
  reg [8-1:0] delete_Key_0_566;
  reg [1-1:0] delete_KeyCompares_0_567;
  reg [3-1:0] delete_KeyCollapse_0_568;
  reg [8-1:0] delete_Data_0_569;
  reg [8-1:0] delete_Key_1_570;
  reg [1-1:0] delete_KeyCompares_1_571;
  reg [3-1:0] delete_KeyCollapse_1_572;
  reg [8-1:0] delete_Data_1_573;
  reg [8-1:0] delete_Key_2_574;
  reg [1-1:0] delete_KeyCompares_2_575;
  reg [3-1:0] delete_KeyCollapse_2_576;
  reg [8-1:0] delete_Data_2_577;
  reg [8-1:0] delete_Key_3_578;
  reg [1-1:0] delete_KeyCompares_3_579;
  reg [3-1:0] delete_KeyCollapse_3_580;
  reg [8-1:0] delete_Data_3_581;
  reg [1-1:0] delete_Found_582;
  reg [8-1:0] delete_Key_583;
  reg [8-1:0] delete_FoundKey_584;
  reg [8-1:0] delete_Data_585;
  reg [6-1:0] delete_BtreeIndex_586;
  reg [3-1:0] delete_StuckIndex_587;
  reg [1-1:0] delete_MergeSuccess_588;
  reg [6-1:0] delete_index_589;
  reg [3-1:0] delete_size_590;
  reg [1-1:0] delete_isLeaf_591;
  reg [6-1:0] delete_nextFree_592;
  reg [8-1:0] delete_Key_0_593;
  reg [1-1:0] delete_KeyCompares_0_594;
  reg [3-1:0] delete_KeyCollapse_0_595;
  reg [8-1:0] delete_Data_0_596;
  reg [8-1:0] delete_Key_1_597;
  reg [1-1:0] delete_KeyCompares_1_598;
  reg [3-1:0] delete_KeyCollapse_1_599;
  reg [8-1:0] delete_Data_1_600;
  reg [8-1:0] delete_Key_2_601;
  reg [1-1:0] delete_KeyCompares_2_602;
  reg [3-1:0] delete_KeyCollapse_2_603;
  reg [8-1:0] delete_Data_2_604;
  reg [8-1:0] delete_Key_3_605;
  reg [1-1:0] delete_KeyCompares_3_606;
  reg [3-1:0] delete_KeyCollapse_3_607;
  reg [8-1:0] delete_Data_3_608;
  reg [1-1:0] delete_Found_609;
  reg [8-1:0] delete_Key_610;
  reg [8-1:0] delete_FoundKey_611;
  reg [8-1:0] delete_Data_612;
  reg [6-1:0] delete_BtreeIndex_613;
  reg [3-1:0] delete_StuckIndex_614;
  reg [1-1:0] delete_MergeSuccess_615;
  reg [8-1:0] delete_childKey_616;
  reg [6-1:0] delete_childData_617;
  reg [6-1:0] delete_indexLeft_618;
  reg [6-1:0] delete_indexRight_619;
  reg [8-1:0] delete_midKey_620;
  reg [1-1:0] delete_success_621;
  reg [1-1:0] delete_test_622;
  reg [6-1:0] delete_next_623;
  reg [6-1:0] delete_root_624;
  reg [1-1:0] delete_isFree_625;
  reg [6-1:0] delete_index_626;
  reg [3-1:0] delete_size_627;
  reg [1-1:0] delete_isLeaf_628;
  reg [6-1:0] delete_nextFree_629;
  reg [8-1:0] delete_Key_0_630;
  reg [1-1:0] delete_KeyCompares_0_631;
  reg [3-1:0] delete_KeyCollapse_0_632;
  reg [8-1:0] delete_Data_0_633;
  reg [8-1:0] delete_Key_1_634;
  reg [1-1:0] delete_KeyCompares_1_635;
  reg [3-1:0] delete_KeyCollapse_1_636;
  reg [8-1:0] delete_Data_1_637;
  reg [8-1:0] delete_Key_2_638;
  reg [1-1:0] delete_KeyCompares_2_639;
  reg [3-1:0] delete_KeyCollapse_2_640;
  reg [8-1:0] delete_Data_2_641;
  reg [8-1:0] delete_Key_3_642;
  reg [1-1:0] delete_KeyCompares_3_643;
  reg [3-1:0] delete_KeyCollapse_3_644;
  reg [8-1:0] delete_Data_3_645;
  reg [1-1:0] delete_Found_646;
  reg [8-1:0] delete_Key_647;
  reg [8-1:0] delete_FoundKey_648;
  reg [8-1:0] delete_Data_649;
  reg [6-1:0] delete_BtreeIndex_650;
  reg [3-1:0] delete_StuckIndex_651;
  reg [1-1:0] delete_MergeSuccess_652;
  reg [6-1:0] delete_index_653;
  reg [3-1:0] delete_size_654;
  reg [1-1:0] delete_isLeaf_655;
  reg [6-1:0] delete_nextFree_656;
  reg [8-1:0] delete_Key_0_657;
  reg [1-1:0] delete_KeyCompares_0_658;
  reg [3-1:0] delete_KeyCollapse_0_659;
  reg [8-1:0] delete_Data_0_660;
  reg [8-1:0] delete_Key_1_661;
  reg [1-1:0] delete_KeyCompares_1_662;
  reg [3-1:0] delete_KeyCollapse_1_663;
  reg [8-1:0] delete_Data_1_664;
  reg [8-1:0] delete_Key_2_665;
  reg [1-1:0] delete_KeyCompares_2_666;
  reg [3-1:0] delete_KeyCollapse_2_667;
  reg [8-1:0] delete_Data_2_668;
  reg [8-1:0] delete_Key_3_669;
  reg [1-1:0] delete_KeyCompares_3_670;
  reg [3-1:0] delete_KeyCollapse_3_671;
  reg [8-1:0] delete_Data_3_672;
  reg [1-1:0] delete_Found_673;
  reg [8-1:0] delete_Key_674;
  reg [8-1:0] delete_FoundKey_675;
  reg [8-1:0] delete_Data_676;
  reg [6-1:0] delete_BtreeIndex_677;
  reg [3-1:0] delete_StuckIndex_678;
  reg [1-1:0] delete_MergeSuccess_679;
  reg [8-1:0] delete_childKey_680;
  reg [3-1:0] delete_leftChild_681;
  reg [3-1:0] delete_rightChild_682;
  reg [6-1:0] delete_childData_683;
  reg [6-1:0] delete_indexLeft_684;
  reg [6-1:0] delete_indexRight_685;
  reg [8-1:0] delete_midKey_686;
  reg [1-1:0] delete_success_687;
  reg [1-1:0] delete_test_688;
  reg [6-1:0] delete_next_689;
  reg [6-1:0] delete_root_690;
  reg [1-1:0] delete_isFree_691;
  reg [6-1:0] delete_index_692;
  reg [3-1:0] delete_size_693;
  reg [1-1:0] delete_isLeaf_694;
  reg [6-1:0] delete_nextFree_695;
  reg [8-1:0] delete_Key_0_696;
  reg [1-1:0] delete_KeyCompares_0_697;
  reg [3-1:0] delete_KeyCollapse_0_698;
  reg [8-1:0] delete_Data_0_699;
  reg [8-1:0] delete_Key_1_700;
  reg [1-1:0] delete_KeyCompares_1_701;
  reg [3-1:0] delete_KeyCollapse_1_702;
  reg [8-1:0] delete_Data_1_703;
  reg [8-1:0] delete_Key_2_704;
  reg [1-1:0] delete_KeyCompares_2_705;
  reg [3-1:0] delete_KeyCollapse_2_706;
  reg [8-1:0] delete_Data_2_707;
  reg [8-1:0] delete_Key_3_708;
  reg [1-1:0] delete_KeyCompares_3_709;
  reg [3-1:0] delete_KeyCollapse_3_710;
  reg [8-1:0] delete_Data_3_711;
  reg [1-1:0] delete_Found_712;
  reg [8-1:0] delete_Key_713;
  reg [8-1:0] delete_FoundKey_714;
  reg [8-1:0] delete_Data_715;
  reg [6-1:0] delete_BtreeIndex_716;
  reg [3-1:0] delete_StuckIndex_717;
  reg [1-1:0] delete_MergeSuccess_718;
  reg [6-1:0] delete_index_719;
  reg [3-1:0] delete_size_720;
  reg [1-1:0] delete_isLeaf_721;
  reg [6-1:0] delete_nextFree_722;
  reg [8-1:0] delete_Key_0_723;
  reg [1-1:0] delete_KeyCompares_0_724;
  reg [3-1:0] delete_KeyCollapse_0_725;
  reg [8-1:0] delete_Data_0_726;
  reg [8-1:0] delete_Key_1_727;
  reg [1-1:0] delete_KeyCompares_1_728;
  reg [3-1:0] delete_KeyCollapse_1_729;
  reg [8-1:0] delete_Data_1_730;
  reg [8-1:0] delete_Key_2_731;
  reg [1-1:0] delete_KeyCompares_2_732;
  reg [3-1:0] delete_KeyCollapse_2_733;
  reg [8-1:0] delete_Data_2_734;
  reg [8-1:0] delete_Key_3_735;
  reg [1-1:0] delete_KeyCompares_3_736;
  reg [3-1:0] delete_KeyCollapse_3_737;
  reg [8-1:0] delete_Data_3_738;
  reg [1-1:0] delete_Found_739;
  reg [8-1:0] delete_Key_740;
  reg [8-1:0] delete_FoundKey_741;
  reg [8-1:0] delete_Data_742;
  reg [6-1:0] delete_BtreeIndex_743;
  reg [3-1:0] delete_StuckIndex_744;
  reg [1-1:0] delete_MergeSuccess_745;
  reg [8-1:0] delete_childKey_746;
  reg [6-1:0] delete_childData_747;
  reg [6-1:0] delete_indexLeft_748;
  reg [6-1:0] delete_indexRight_749;
  reg [8-1:0] delete_midKey_750;
  reg [1-1:0] delete_success_751;
  reg [1-1:0] delete_test_752;
  reg [6-1:0] delete_next_753;
  reg [6-1:0] delete_root_754;
  reg [1-1:0] delete_isFree_755;
  reg [6-1:0] delete_index_756;
  reg [3-1:0] delete_size_757;
  reg [1-1:0] delete_isLeaf_758;
  reg [6-1:0] delete_nextFree_759;
  reg [8-1:0] delete_Key_0_760;
  reg [1-1:0] delete_KeyCompares_0_761;
  reg [3-1:0] delete_KeyCollapse_0_762;
  reg [8-1:0] delete_Data_0_763;
  reg [8-1:0] delete_Key_1_764;
  reg [1-1:0] delete_KeyCompares_1_765;
  reg [3-1:0] delete_KeyCollapse_1_766;
  reg [8-1:0] delete_Data_1_767;
  reg [8-1:0] delete_Key_2_768;
  reg [1-1:0] delete_KeyCompares_2_769;
  reg [3-1:0] delete_KeyCollapse_2_770;
  reg [8-1:0] delete_Data_2_771;
  reg [8-1:0] delete_Key_3_772;
  reg [1-1:0] delete_KeyCompares_3_773;
  reg [3-1:0] delete_KeyCollapse_3_774;
  reg [8-1:0] delete_Data_3_775;
  reg [1-1:0] delete_Found_776;
  reg [8-1:0] delete_Key_777;
  reg [8-1:0] delete_FoundKey_778;
  reg [8-1:0] delete_Data_779;
  reg [6-1:0] delete_BtreeIndex_780;
  reg [3-1:0] delete_StuckIndex_781;
  reg [1-1:0] delete_MergeSuccess_782;
  reg [6-1:0] delete_index_783;
  reg [3-1:0] delete_size_784;
  reg [1-1:0] delete_isLeaf_785;
  reg [6-1:0] delete_nextFree_786;
  reg [8-1:0] delete_Key_0_787;
  reg [1-1:0] delete_KeyCompares_0_788;
  reg [3-1:0] delete_KeyCollapse_0_789;
  reg [8-1:0] delete_Data_0_790;
  reg [8-1:0] delete_Key_1_791;
  reg [1-1:0] delete_KeyCompares_1_792;
  reg [3-1:0] delete_KeyCollapse_1_793;
  reg [8-1:0] delete_Data_1_794;
  reg [8-1:0] delete_Key_2_795;
  reg [1-1:0] delete_KeyCompares_2_796;
  reg [3-1:0] delete_KeyCollapse_2_797;
  reg [8-1:0] delete_Data_2_798;
  reg [8-1:0] delete_Key_3_799;
  reg [1-1:0] delete_KeyCompares_3_800;
  reg [3-1:0] delete_KeyCollapse_3_801;
  reg [8-1:0] delete_Data_3_802;
  reg [1-1:0] delete_Found_803;
  reg [8-1:0] delete_Key_804;
  reg [8-1:0] delete_FoundKey_805;
  reg [8-1:0] delete_Data_806;
  reg [6-1:0] delete_BtreeIndex_807;
  reg [3-1:0] delete_StuckIndex_808;
  reg [1-1:0] delete_MergeSuccess_809;
  reg [8-1:0] delete_childKey_810;
  reg [3-1:0] delete_leftChild_811;
  reg [3-1:0] delete_rightChild_812;
  reg [6-1:0] delete_childData_813;
  reg [6-1:0] delete_indexLeft_814;
  reg [6-1:0] delete_indexRight_815;
  reg [8-1:0] delete_midKey_816;
  reg [1-1:0] delete_success_817;
  reg [1-1:0] delete_test_818;
  reg [6-1:0] delete_next_819;
  reg [6-1:0] delete_root_820;
  reg [1-1:0] delete_isFree_821;
  reg [6-1:0] delete_index_822;
  reg [3-1:0] delete_size_823;
  reg [1-1:0] delete_isLeaf_824;
  reg [6-1:0] delete_nextFree_825;
  reg [8-1:0] delete_Key_0_826;
  reg [1-1:0] delete_KeyCompares_0_827;
  reg [3-1:0] delete_KeyCollapse_0_828;
  reg [8-1:0] delete_Data_0_829;
  reg [8-1:0] delete_Key_1_830;
  reg [1-1:0] delete_KeyCompares_1_831;
  reg [3-1:0] delete_KeyCollapse_1_832;
  reg [8-1:0] delete_Data_1_833;
  reg [8-1:0] delete_Key_2_834;
  reg [1-1:0] delete_KeyCompares_2_835;
  reg [3-1:0] delete_KeyCollapse_2_836;
  reg [8-1:0] delete_Data_2_837;
  reg [8-1:0] delete_Key_3_838;
  reg [1-1:0] delete_KeyCompares_3_839;
  reg [3-1:0] delete_KeyCollapse_3_840;
  reg [8-1:0] delete_Data_3_841;
  reg [1-1:0] delete_Found_842;
  reg [8-1:0] delete_Key_843;
  reg [8-1:0] delete_FoundKey_844;
  reg [8-1:0] delete_Data_845;
  reg [6-1:0] delete_BtreeIndex_846;
  reg [3-1:0] delete_StuckIndex_847;
  reg [1-1:0] delete_MergeSuccess_848;
  reg [6-1:0] delete_index_849;
  reg [3-1:0] delete_size_850;
  reg [1-1:0] delete_isLeaf_851;
  reg [6-1:0] delete_nextFree_852;
  reg [8-1:0] delete_Key_0_853;
  reg [1-1:0] delete_KeyCompares_0_854;
  reg [3-1:0] delete_KeyCollapse_0_855;
  reg [8-1:0] delete_Data_0_856;
  reg [8-1:0] delete_Key_1_857;
  reg [1-1:0] delete_KeyCompares_1_858;
  reg [3-1:0] delete_KeyCollapse_1_859;
  reg [8-1:0] delete_Data_1_860;
  reg [8-1:0] delete_Key_2_861;
  reg [1-1:0] delete_KeyCompares_2_862;
  reg [3-1:0] delete_KeyCollapse_2_863;
  reg [8-1:0] delete_Data_2_864;
  reg [8-1:0] delete_Key_3_865;
  reg [1-1:0] delete_KeyCompares_3_866;
  reg [3-1:0] delete_KeyCollapse_3_867;
  reg [8-1:0] delete_Data_3_868;
  reg [1-1:0] delete_Found_869;
  reg [8-1:0] delete_Key_870;
  reg [8-1:0] delete_FoundKey_871;
  reg [8-1:0] delete_Data_872;
  reg [6-1:0] delete_BtreeIndex_873;
  reg [3-1:0] delete_StuckIndex_874;
  reg [1-1:0] delete_MergeSuccess_875;
  reg [8-1:0] delete_childKey_876;
  reg [6-1:0] delete_childData_877;
  reg [6-1:0] delete_indexLeft_878;
  reg [6-1:0] delete_indexRight_879;
  reg [8-1:0] delete_midKey_880;
  reg [1-1:0] delete_success_881;
  reg [1-1:0] delete_test_882;
  reg [6-1:0] delete_next_883;
  reg [6-1:0] delete_root_884;
  reg [1-1:0] delete_isFree_885;
  reg [6-1:0] delete_index_886;
  reg [3-1:0] delete_size_887;
  reg [1-1:0] delete_isLeaf_888;
  reg [6-1:0] delete_nextFree_889;
  reg [8-1:0] delete_Key_0_890;
  reg [1-1:0] delete_KeyCompares_0_891;
  reg [3-1:0] delete_KeyCollapse_0_892;
  reg [8-1:0] delete_Data_0_893;
  reg [8-1:0] delete_Key_1_894;
  reg [1-1:0] delete_KeyCompares_1_895;
  reg [3-1:0] delete_KeyCollapse_1_896;
  reg [8-1:0] delete_Data_1_897;
  reg [8-1:0] delete_Key_2_898;
  reg [1-1:0] delete_KeyCompares_2_899;
  reg [3-1:0] delete_KeyCollapse_2_900;
  reg [8-1:0] delete_Data_2_901;
  reg [8-1:0] delete_Key_3_902;
  reg [1-1:0] delete_KeyCompares_3_903;
  reg [3-1:0] delete_KeyCollapse_3_904;
  reg [8-1:0] delete_Data_3_905;
  reg [1-1:0] delete_Found_906;
  reg [8-1:0] delete_Key_907;
  reg [8-1:0] delete_FoundKey_908;
  reg [8-1:0] delete_Data_909;
  reg [6-1:0] delete_BtreeIndex_910;
  reg [3-1:0] delete_StuckIndex_911;
  reg [1-1:0] delete_MergeSuccess_912;
  reg [6-1:0] delete_index_913;
  reg [3-1:0] delete_size_914;
  reg [1-1:0] delete_isLeaf_915;
  reg [6-1:0] delete_nextFree_916;
  reg [8-1:0] delete_Key_0_917;
  reg [1-1:0] delete_KeyCompares_0_918;
  reg [3-1:0] delete_KeyCollapse_0_919;
  reg [8-1:0] delete_Data_0_920;
  reg [8-1:0] delete_Key_1_921;
  reg [1-1:0] delete_KeyCompares_1_922;
  reg [3-1:0] delete_KeyCollapse_1_923;
  reg [8-1:0] delete_Data_1_924;
  reg [8-1:0] delete_Key_2_925;
  reg [1-1:0] delete_KeyCompares_2_926;
  reg [3-1:0] delete_KeyCollapse_2_927;
  reg [8-1:0] delete_Data_2_928;
  reg [8-1:0] delete_Key_3_929;
  reg [1-1:0] delete_KeyCompares_3_930;
  reg [3-1:0] delete_KeyCollapse_3_931;
  reg [8-1:0] delete_Data_3_932;
  reg [1-1:0] delete_Found_933;
  reg [8-1:0] delete_Key_934;
  reg [8-1:0] delete_FoundKey_935;
  reg [8-1:0] delete_Data_936;
  reg [6-1:0] delete_BtreeIndex_937;
  reg [3-1:0] delete_StuckIndex_938;
  reg [1-1:0] delete_MergeSuccess_939;
  reg [8-1:0] delete_childKey_940;
  reg [3-1:0] delete_leftChild_941;
  reg [3-1:0] delete_rightChild_942;
  reg [6-1:0] delete_childData_943;
  reg [6-1:0] delete_indexLeft_944;
  reg [6-1:0] delete_indexRight_945;
  reg [8-1:0] delete_midKey_946;
  reg [1-1:0] delete_success_947;
  reg [1-1:0] delete_test_948;
  reg [6-1:0] delete_next_949;
  reg [6-1:0] delete_root_950;
  reg [1-1:0] delete_isFree_951;
  reg [6-1:0] delete_index_952;
  reg [3-1:0] delete_size_953;
  reg [1-1:0] delete_isLeaf_954;
  reg [6-1:0] delete_nextFree_955;
  reg [8-1:0] delete_Key_0_956;
  reg [1-1:0] delete_KeyCompares_0_957;
  reg [3-1:0] delete_KeyCollapse_0_958;
  reg [8-1:0] delete_Data_0_959;
  reg [8-1:0] delete_Key_1_960;
  reg [1-1:0] delete_KeyCompares_1_961;
  reg [3-1:0] delete_KeyCollapse_1_962;
  reg [8-1:0] delete_Data_1_963;
  reg [8-1:0] delete_Key_2_964;
  reg [1-1:0] delete_KeyCompares_2_965;
  reg [3-1:0] delete_KeyCollapse_2_966;
  reg [8-1:0] delete_Data_2_967;
  reg [8-1:0] delete_Key_3_968;
  reg [1-1:0] delete_KeyCompares_3_969;
  reg [3-1:0] delete_KeyCollapse_3_970;
  reg [8-1:0] delete_Data_3_971;
  reg [1-1:0] delete_Found_972;
  reg [8-1:0] delete_Key_973;
  reg [8-1:0] delete_FoundKey_974;
  reg [8-1:0] delete_Data_975;
  reg [6-1:0] delete_BtreeIndex_976;
  reg [3-1:0] delete_StuckIndex_977;
  reg [1-1:0] delete_MergeSuccess_978;
  reg [6-1:0] delete_index_979;
  reg [3-1:0] delete_size_980;
  reg [1-1:0] delete_isLeaf_981;
  reg [6-1:0] delete_nextFree_982;
  reg [8-1:0] delete_Key_0_983;
  reg [1-1:0] delete_KeyCompares_0_984;
  reg [3-1:0] delete_KeyCollapse_0_985;
  reg [8-1:0] delete_Data_0_986;
  reg [8-1:0] delete_Key_1_987;
  reg [1-1:0] delete_KeyCompares_1_988;
  reg [3-1:0] delete_KeyCollapse_1_989;
  reg [8-1:0] delete_Data_1_990;
  reg [8-1:0] delete_Key_2_991;
  reg [1-1:0] delete_KeyCompares_2_992;
  reg [3-1:0] delete_KeyCollapse_2_993;
  reg [8-1:0] delete_Data_2_994;
  reg [8-1:0] delete_Key_3_995;
  reg [1-1:0] delete_KeyCompares_3_996;
  reg [3-1:0] delete_KeyCollapse_3_997;
  reg [8-1:0] delete_Data_3_998;
  reg [1-1:0] delete_Found_999;
  reg [8-1:0] delete_Key_1000;
  reg [8-1:0] delete_FoundKey_1001;
  reg [8-1:0] delete_Data_1002;
  reg [6-1:0] delete_BtreeIndex_1003;
  reg [3-1:0] delete_StuckIndex_1004;
  reg [1-1:0] delete_MergeSuccess_1005;
  reg [8-1:0] delete_childKey_1006;
  reg [6-1:0] delete_childData_1007;
  reg [6-1:0] delete_indexLeft_1008;
  reg [6-1:0] delete_indexRight_1009;
  reg [8-1:0] delete_midKey_1010;
  reg [1-1:0] delete_success_1011;
  reg [1-1:0] delete_test_1012;
  reg [6-1:0] delete_next_1013;
  reg [6-1:0] delete_root_1014;
  reg [1-1:0] delete_isFree_1015;
  reg [6-1:0] delete_index_1016;
  reg [3-1:0] delete_size_1017;
  reg [1-1:0] delete_isLeaf_1018;
  reg [6-1:0] delete_nextFree_1019;
  reg [8-1:0] delete_Key_0_1020;
  reg [1-1:0] delete_KeyCompares_0_1021;
  reg [3-1:0] delete_KeyCollapse_0_1022;
  reg [8-1:0] delete_Data_0_1023;
  reg [8-1:0] delete_Key_1_1024;
  reg [1-1:0] delete_KeyCompares_1_1025;
  reg [3-1:0] delete_KeyCollapse_1_1026;
  reg [8-1:0] delete_Data_1_1027;
  reg [8-1:0] delete_Key_2_1028;
  reg [1-1:0] delete_KeyCompares_2_1029;
  reg [3-1:0] delete_KeyCollapse_2_1030;
  reg [8-1:0] delete_Data_2_1031;
  reg [8-1:0] delete_Key_3_1032;
  reg [1-1:0] delete_KeyCompares_3_1033;
  reg [3-1:0] delete_KeyCollapse_3_1034;
  reg [8-1:0] delete_Data_3_1035;
  reg [1-1:0] delete_Found_1036;
  reg [8-1:0] delete_Key_1037;
  reg [8-1:0] delete_FoundKey_1038;
  reg [8-1:0] delete_Data_1039;
  reg [6-1:0] delete_BtreeIndex_1040;
  reg [3-1:0] delete_StuckIndex_1041;
  reg [1-1:0] delete_MergeSuccess_1042;
  reg [6-1:0] delete_index_1043;
  reg [3-1:0] delete_size_1044;
  reg [1-1:0] delete_isLeaf_1045;
  reg [6-1:0] delete_nextFree_1046;
  reg [8-1:0] delete_Key_0_1047;
  reg [1-1:0] delete_KeyCompares_0_1048;
  reg [3-1:0] delete_KeyCollapse_0_1049;
  reg [8-1:0] delete_Data_0_1050;
  reg [8-1:0] delete_Key_1_1051;
  reg [1-1:0] delete_KeyCompares_1_1052;
  reg [3-1:0] delete_KeyCollapse_1_1053;
  reg [8-1:0] delete_Data_1_1054;
  reg [8-1:0] delete_Key_2_1055;
  reg [1-1:0] delete_KeyCompares_2_1056;
  reg [3-1:0] delete_KeyCollapse_2_1057;
  reg [8-1:0] delete_Data_2_1058;
  reg [8-1:0] delete_Key_3_1059;
  reg [1-1:0] delete_KeyCompares_3_1060;
  reg [3-1:0] delete_KeyCollapse_3_1061;
  reg [8-1:0] delete_Data_3_1062;
  reg [1-1:0] delete_Found_1063;
  reg [8-1:0] delete_Key_1064;
  reg [8-1:0] delete_FoundKey_1065;
  reg [8-1:0] delete_Data_1066;
  reg [6-1:0] delete_BtreeIndex_1067;
  reg [3-1:0] delete_StuckIndex_1068;
  reg [1-1:0] delete_MergeSuccess_1069;
  reg [8-1:0] delete_childKey_1070;
  reg [3-1:0] delete_leftChild_1071;
  reg [3-1:0] delete_rightChild_1072;
  reg [6-1:0] delete_childData_1073;
  reg [6-1:0] delete_indexLeft_1074;
  reg [6-1:0] delete_indexRight_1075;
  reg [8-1:0] delete_midKey_1076;
  reg [1-1:0] delete_success_1077;
  reg [1-1:0] delete_test_1078;
  reg [6-1:0] delete_next_1079;
  reg [6-1:0] delete_root_1080;
  reg [1-1:0] delete_isFree_1081;
  reg [6-1:0] delete_index_1082;
  reg [3-1:0] delete_size_1083;
  reg [1-1:0] delete_isLeaf_1084;
  reg [6-1:0] delete_nextFree_1085;
  reg [8-1:0] delete_Key_0_1086;
  reg [1-1:0] delete_KeyCompares_0_1087;
  reg [3-1:0] delete_KeyCollapse_0_1088;
  reg [8-1:0] delete_Data_0_1089;
  reg [8-1:0] delete_Key_1_1090;
  reg [1-1:0] delete_KeyCompares_1_1091;
  reg [3-1:0] delete_KeyCollapse_1_1092;
  reg [8-1:0] delete_Data_1_1093;
  reg [8-1:0] delete_Key_2_1094;
  reg [1-1:0] delete_KeyCompares_2_1095;
  reg [3-1:0] delete_KeyCollapse_2_1096;
  reg [8-1:0] delete_Data_2_1097;
  reg [8-1:0] delete_Key_3_1098;
  reg [1-1:0] delete_KeyCompares_3_1099;
  reg [3-1:0] delete_KeyCollapse_3_1100;
  reg [8-1:0] delete_Data_3_1101;
  reg [1-1:0] delete_Found_1102;
  reg [8-1:0] delete_Key_1103;
  reg [8-1:0] delete_FoundKey_1104;
  reg [8-1:0] delete_Data_1105;
  reg [6-1:0] delete_BtreeIndex_1106;
  reg [3-1:0] delete_StuckIndex_1107;
  reg [1-1:0] delete_MergeSuccess_1108;
  reg [6-1:0] delete_index_1109;
  reg [3-1:0] delete_size_1110;
  reg [1-1:0] delete_isLeaf_1111;
  reg [6-1:0] delete_nextFree_1112;
  reg [8-1:0] delete_Key_0_1113;
  reg [1-1:0] delete_KeyCompares_0_1114;
  reg [3-1:0] delete_KeyCollapse_0_1115;
  reg [8-1:0] delete_Data_0_1116;
  reg [8-1:0] delete_Key_1_1117;
  reg [1-1:0] delete_KeyCompares_1_1118;
  reg [3-1:0] delete_KeyCollapse_1_1119;
  reg [8-1:0] delete_Data_1_1120;
  reg [8-1:0] delete_Key_2_1121;
  reg [1-1:0] delete_KeyCompares_2_1122;
  reg [3-1:0] delete_KeyCollapse_2_1123;
  reg [8-1:0] delete_Data_2_1124;
  reg [8-1:0] delete_Key_3_1125;
  reg [1-1:0] delete_KeyCompares_3_1126;
  reg [3-1:0] delete_KeyCollapse_3_1127;
  reg [8-1:0] delete_Data_3_1128;
  reg [1-1:0] delete_Found_1129;
  reg [8-1:0] delete_Key_1130;
  reg [8-1:0] delete_FoundKey_1131;
  reg [8-1:0] delete_Data_1132;
  reg [6-1:0] delete_BtreeIndex_1133;
  reg [3-1:0] delete_StuckIndex_1134;
  reg [1-1:0] delete_MergeSuccess_1135;
  reg [8-1:0] delete_childKey_1136;
  reg [6-1:0] delete_childData_1137;
  reg [6-1:0] delete_indexLeft_1138;
  reg [6-1:0] delete_indexRight_1139;
  reg [8-1:0] delete_midKey_1140;
  reg [1-1:0] delete_success_1141;
  reg [1-1:0] delete_test_1142;
  reg [6-1:0] delete_next_1143;
  reg [6-1:0] delete_root_1144;
  reg [1-1:0] delete_isFree_1145;
  reg [6-1:0] delete_index_1146;
  reg [3-1:0] delete_size_1147;
  reg [1-1:0] delete_isLeaf_1148;
  reg [6-1:0] delete_nextFree_1149;
  reg [8-1:0] delete_Key_0_1150;
  reg [1-1:0] delete_KeyCompares_0_1151;
  reg [3-1:0] delete_KeyCollapse_0_1152;
  reg [8-1:0] delete_Data_0_1153;
  reg [8-1:0] delete_Key_1_1154;
  reg [1-1:0] delete_KeyCompares_1_1155;
  reg [3-1:0] delete_KeyCollapse_1_1156;
  reg [8-1:0] delete_Data_1_1157;
  reg [8-1:0] delete_Key_2_1158;
  reg [1-1:0] delete_KeyCompares_2_1159;
  reg [3-1:0] delete_KeyCollapse_2_1160;
  reg [8-1:0] delete_Data_2_1161;
  reg [8-1:0] delete_Key_3_1162;
  reg [1-1:0] delete_KeyCompares_3_1163;
  reg [3-1:0] delete_KeyCollapse_3_1164;
  reg [8-1:0] delete_Data_3_1165;
  reg [1-1:0] delete_Found_1166;
  reg [8-1:0] delete_Key_1167;
  reg [8-1:0] delete_FoundKey_1168;
  reg [8-1:0] delete_Data_1169;
  reg [6-1:0] delete_BtreeIndex_1170;
  reg [3-1:0] delete_StuckIndex_1171;
  reg [1-1:0] delete_MergeSuccess_1172;
  reg [6-1:0] delete_index_1173;
  reg [3-1:0] delete_size_1174;
  reg [1-1:0] delete_isLeaf_1175;
  reg [6-1:0] delete_nextFree_1176;
  reg [8-1:0] delete_Key_0_1177;
  reg [1-1:0] delete_KeyCompares_0_1178;
  reg [3-1:0] delete_KeyCollapse_0_1179;
  reg [8-1:0] delete_Data_0_1180;
  reg [8-1:0] delete_Key_1_1181;
  reg [1-1:0] delete_KeyCompares_1_1182;
  reg [3-1:0] delete_KeyCollapse_1_1183;
  reg [8-1:0] delete_Data_1_1184;
  reg [8-1:0] delete_Key_2_1185;
  reg [1-1:0] delete_KeyCompares_2_1186;
  reg [3-1:0] delete_KeyCollapse_2_1187;
  reg [8-1:0] delete_Data_2_1188;
  reg [8-1:0] delete_Key_3_1189;
  reg [1-1:0] delete_KeyCompares_3_1190;
  reg [3-1:0] delete_KeyCollapse_3_1191;
  reg [8-1:0] delete_Data_3_1192;
  reg [1-1:0] delete_Found_1193;
  reg [8-1:0] delete_Key_1194;
  reg [8-1:0] delete_FoundKey_1195;
  reg [8-1:0] delete_Data_1196;
  reg [6-1:0] delete_BtreeIndex_1197;
  reg [3-1:0] delete_StuckIndex_1198;
  reg [1-1:0] delete_MergeSuccess_1199;
  reg [8-1:0] delete_childKey_1200;
  reg [3-1:0] delete_leftChild_1201;
  reg [3-1:0] delete_rightChild_1202;
  reg [6-1:0] delete_childData_1203;
  reg [6-1:0] delete_indexLeft_1204;
  reg [6-1:0] delete_indexRight_1205;
  reg [8-1:0] delete_midKey_1206;
  reg [1-1:0] delete_success_1207;
  reg [1-1:0] delete_test_1208;
  reg [6-1:0] delete_next_1209;
  reg [6-1:0] delete_root_1210;
  reg [1-1:0] delete_isFree_1211;
  integer delete_pc;
  integer delete_stop;
  integer delete_returnCode;
  integer delete_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      delete_pc <= 0;
      delete_stop <= 0;
      delete_returnCode <= 0;
      delete_index_0 <= 0;
      delete_size_1 <= 0;
      delete_isLeaf_2 <= 0;
      delete_nextFree_3 <= 0;
      delete_Key_0_4 <= 0;
      delete_KeyCompares_0_5 <= 0;
      delete_KeyCollapse_0_6 <= 0;
      delete_Data_0_7 <= 0;
      delete_Key_1_8 <= 0;
      delete_KeyCompares_1_9 <= 0;
      delete_KeyCollapse_1_10 <= 0;
      delete_Data_1_11 <= 0;
      delete_Key_2_12 <= 0;
      delete_KeyCompares_2_13 <= 0;
      delete_KeyCollapse_2_14 <= 0;
      delete_Data_2_15 <= 0;
      delete_Key_3_16 <= 0;
      delete_KeyCompares_3_17 <= 0;
      delete_KeyCollapse_3_18 <= 0;
      delete_Data_3_19 <= 0;
      delete_stuckKeys_1_index_20 <= 0;
      delete_stuckKeys_2_index_21 <= 0;
      delete_stuckKeys_2_value_22 <= 0;
      delete_stuckKeys_2_value_23 <= 0;
      delete_stuckKeys_2_value_24 <= 0;
      delete_stuckKeys_2_value_25 <= 0;
      delete_stuckData_3_index_26 <= 0;
      delete_stuckData_4_index_27 <= 0;
      delete_stuckData_4_value_28 <= 0;
      delete_stuckData_4_value_29 <= 0;
      delete_stuckData_4_value_30 <= 0;
      delete_stuckData_4_value_31 <= 0;
      delete_stuckSize_5_index_32 <= 0;
      delete_stuckSize_6_index_33 <= 0;
      delete_stuckSize_6_value_34 <= 0;
      delete_stuckIsLeaf_7_index_35 <= 0;
      delete_stuckIsLeaf_8_index_36 <= 0;
      delete_stuckIsLeaf_8_value_37 <= 0;
      delete_Found_38 <= 0;
      delete_Key_39 <= 0;
      delete_FoundKey_40 <= 0;
      delete_Data_41 <= 0;
      delete_BtreeIndex_42 <= 0;
      delete_StuckIndex_43 <= 0;
      delete_MergeSuccess_44 <= 0;
      delete_i_45 <= 0;
      delete_k_46 <= 0;
      delete_l_47 <= 0;
      delete_index_48 <= 0;
      delete_size_49 <= 0;
      delete_isLeaf_50 <= 0;
      delete_nextFree_51 <= 0;
      delete_Key_0_52 <= 0;
      delete_KeyCompares_0_53 <= 0;
      delete_KeyCollapse_0_54 <= 0;
      delete_Data_0_55 <= 0;
      delete_Key_1_56 <= 0;
      delete_KeyCompares_1_57 <= 0;
      delete_KeyCollapse_1_58 <= 0;
      delete_Data_1_59 <= 0;
      delete_Key_2_60 <= 0;
      delete_KeyCompares_2_61 <= 0;
      delete_KeyCollapse_2_62 <= 0;
      delete_Data_2_63 <= 0;
      delete_Key_3_64 <= 0;
      delete_KeyCompares_3_65 <= 0;
      delete_KeyCollapse_3_66 <= 0;
      delete_Data_3_67 <= 0;
      delete_Found_68 <= 0;
      delete_Key_69 <= 0;
      delete_FoundKey_70 <= 0;
      delete_Data_71 <= 0;
      delete_BtreeIndex_72 <= 0;
      delete_StuckIndex_73 <= 0;
      delete_MergeSuccess_74 <= 0;
      delete_index_75 <= 0;
      delete_size_76 <= 0;
      delete_isLeaf_77 <= 0;
      delete_nextFree_78 <= 0;
      delete_Key_0_79 <= 0;
      delete_KeyCompares_0_80 <= 0;
      delete_KeyCollapse_0_81 <= 0;
      delete_Data_0_82 <= 0;
      delete_Key_1_83 <= 0;
      delete_KeyCompares_1_84 <= 0;
      delete_KeyCollapse_1_85 <= 0;
      delete_Data_1_86 <= 0;
      delete_Key_2_87 <= 0;
      delete_KeyCompares_2_88 <= 0;
      delete_KeyCollapse_2_89 <= 0;
      delete_Data_2_90 <= 0;
      delete_Key_3_91 <= 0;
      delete_KeyCompares_3_92 <= 0;
      delete_KeyCollapse_3_93 <= 0;
      delete_Data_3_94 <= 0;
      delete_Found_95 <= 0;
      delete_Key_96 <= 0;
      delete_FoundKey_97 <= 0;
      delete_Data_98 <= 0;
      delete_BtreeIndex_99 <= 0;
      delete_StuckIndex_100 <= 0;
      delete_MergeSuccess_101 <= 0;
      delete_position_102 <= 0;
      delete_index_103 <= 0;
      delete_index1_104 <= 0;
      delete_within_105 <= 0;
      delete_isLeaf_106 <= 0;
      delete_index_107 <= 0;
      delete_size_108 <= 0;
      delete_isLeaf_109 <= 0;
      delete_nextFree_110 <= 0;
      delete_Key_0_111 <= 0;
      delete_KeyCompares_0_112 <= 0;
      delete_KeyCollapse_0_113 <= 0;
      delete_Data_0_114 <= 0;
      delete_Key_1_115 <= 0;
      delete_KeyCompares_1_116 <= 0;
      delete_KeyCollapse_1_117 <= 0;
      delete_Data_1_118 <= 0;
      delete_Key_2_119 <= 0;
      delete_KeyCompares_2_120 <= 0;
      delete_KeyCollapse_2_121 <= 0;
      delete_Data_2_122 <= 0;
      delete_Key_3_123 <= 0;
      delete_KeyCompares_3_124 <= 0;
      delete_KeyCollapse_3_125 <= 0;
      delete_Data_3_126 <= 0;
      delete_Found_127 <= 0;
      delete_Key_128 <= 0;
      delete_FoundKey_129 <= 0;
      delete_Data_130 <= 0;
      delete_BtreeIndex_131 <= 0;
      delete_StuckIndex_132 <= 0;
      delete_MergeSuccess_133 <= 0;
      delete_index_134 <= 0;
      delete_size_135 <= 0;
      delete_isLeaf_136 <= 0;
      delete_nextFree_137 <= 0;
      delete_Key_0_138 <= 0;
      delete_KeyCompares_0_139 <= 0;
      delete_KeyCollapse_0_140 <= 0;
      delete_Data_0_141 <= 0;
      delete_Key_1_142 <= 0;
      delete_KeyCompares_1_143 <= 0;
      delete_KeyCollapse_1_144 <= 0;
      delete_Data_1_145 <= 0;
      delete_Key_2_146 <= 0;
      delete_KeyCompares_2_147 <= 0;
      delete_KeyCollapse_2_148 <= 0;
      delete_Data_2_149 <= 0;
      delete_Key_3_150 <= 0;
      delete_KeyCompares_3_151 <= 0;
      delete_KeyCollapse_3_152 <= 0;
      delete_Data_3_153 <= 0;
      delete_Found_154 <= 0;
      delete_Key_155 <= 0;
      delete_FoundKey_156 <= 0;
      delete_Data_157 <= 0;
      delete_BtreeIndex_158 <= 0;
      delete_StuckIndex_159 <= 0;
      delete_MergeSuccess_160 <= 0;
      delete_index_161 <= 0;
      delete_size_162 <= 0;
      delete_isLeaf_163 <= 0;
      delete_nextFree_164 <= 0;
      delete_Key_0_165 <= 0;
      delete_KeyCompares_0_166 <= 0;
      delete_KeyCollapse_0_167 <= 0;
      delete_Data_0_168 <= 0;
      delete_Key_1_169 <= 0;
      delete_KeyCompares_1_170 <= 0;
      delete_KeyCollapse_1_171 <= 0;
      delete_Data_1_172 <= 0;
      delete_Key_2_173 <= 0;
      delete_KeyCompares_2_174 <= 0;
      delete_KeyCollapse_2_175 <= 0;
      delete_Data_2_176 <= 0;
      delete_Key_3_177 <= 0;
      delete_KeyCompares_3_178 <= 0;
      delete_KeyCollapse_3_179 <= 0;
      delete_Data_3_180 <= 0;
      delete_Found_181 <= 0;
      delete_Key_182 <= 0;
      delete_FoundKey_183 <= 0;
      delete_Data_184 <= 0;
      delete_BtreeIndex_185 <= 0;
      delete_StuckIndex_186 <= 0;
      delete_MergeSuccess_187 <= 0;
      delete_childKey_188 <= 0;
      delete_childData_189 <= 0;
      delete_indexLeft_190 <= 0;
      delete_indexRight_191 <= 0;
      delete_midKey_192 <= 0;
      delete_success_193 <= 0;
      delete_test_194 <= 0;
      delete_next_195 <= 0;
      delete_freeNext_9_index_196 <= 0;
      delete_freeNext_10_index_197 <= 0;
      delete_freeNext_10_value_198 <= 0;
      delete_stuckIsFree_11_index_199 <= 0;
      delete_stuckIsFree_11_value_200 <= 0;
      delete_root_201 <= 0;
      delete_isFree_202 <= 0;
      delete_next_203 <= 0;
      delete_root_204 <= 0;
      delete_isFree_205 <= 0;
      delete_index_206 <= 0;
      delete_size_207 <= 0;
      delete_isLeaf_208 <= 0;
      delete_nextFree_209 <= 0;
      delete_Key_0_210 <= 0;
      delete_KeyCompares_0_211 <= 0;
      delete_KeyCollapse_0_212 <= 0;
      delete_Data_0_213 <= 0;
      delete_Key_1_214 <= 0;
      delete_KeyCompares_1_215 <= 0;
      delete_KeyCollapse_1_216 <= 0;
      delete_Data_1_217 <= 0;
      delete_Key_2_218 <= 0;
      delete_KeyCompares_2_219 <= 0;
      delete_KeyCollapse_2_220 <= 0;
      delete_Data_2_221 <= 0;
      delete_Key_3_222 <= 0;
      delete_KeyCompares_3_223 <= 0;
      delete_KeyCollapse_3_224 <= 0;
      delete_Data_3_225 <= 0;
      delete_Found_226 <= 0;
      delete_Key_227 <= 0;
      delete_FoundKey_228 <= 0;
      delete_Data_229 <= 0;
      delete_BtreeIndex_230 <= 0;
      delete_StuckIndex_231 <= 0;
      delete_MergeSuccess_232 <= 0;
      delete_index_233 <= 0;
      delete_size_234 <= 0;
      delete_isLeaf_235 <= 0;
      delete_nextFree_236 <= 0;
      delete_Key_0_237 <= 0;
      delete_KeyCompares_0_238 <= 0;
      delete_KeyCollapse_0_239 <= 0;
      delete_Data_0_240 <= 0;
      delete_Key_1_241 <= 0;
      delete_KeyCompares_1_242 <= 0;
      delete_KeyCollapse_1_243 <= 0;
      delete_Data_1_244 <= 0;
      delete_Key_2_245 <= 0;
      delete_KeyCompares_2_246 <= 0;
      delete_KeyCollapse_2_247 <= 0;
      delete_Data_2_248 <= 0;
      delete_Key_3_249 <= 0;
      delete_KeyCompares_3_250 <= 0;
      delete_KeyCollapse_3_251 <= 0;
      delete_Data_3_252 <= 0;
      delete_Found_253 <= 0;
      delete_Key_254 <= 0;
      delete_FoundKey_255 <= 0;
      delete_Data_256 <= 0;
      delete_BtreeIndex_257 <= 0;
      delete_StuckIndex_258 <= 0;
      delete_MergeSuccess_259 <= 0;
      delete_index_260 <= 0;
      delete_size_261 <= 0;
      delete_isLeaf_262 <= 0;
      delete_nextFree_263 <= 0;
      delete_Key_0_264 <= 0;
      delete_KeyCompares_0_265 <= 0;
      delete_KeyCollapse_0_266 <= 0;
      delete_Data_0_267 <= 0;
      delete_Key_1_268 <= 0;
      delete_KeyCompares_1_269 <= 0;
      delete_KeyCollapse_1_270 <= 0;
      delete_Data_1_271 <= 0;
      delete_Key_2_272 <= 0;
      delete_KeyCompares_2_273 <= 0;
      delete_KeyCollapse_2_274 <= 0;
      delete_Data_2_275 <= 0;
      delete_Key_3_276 <= 0;
      delete_KeyCompares_3_277 <= 0;
      delete_KeyCollapse_3_278 <= 0;
      delete_Data_3_279 <= 0;
      delete_Found_280 <= 0;
      delete_Key_281 <= 0;
      delete_FoundKey_282 <= 0;
      delete_Data_283 <= 0;
      delete_BtreeIndex_284 <= 0;
      delete_StuckIndex_285 <= 0;
      delete_MergeSuccess_286 <= 0;
      delete_childKey_287 <= 0;
      delete_leftChild_288 <= 0;
      delete_rightChild_289 <= 0;
      delete_childData_290 <= 0;
      delete_indexLeft_291 <= 0;
      delete_indexRight_292 <= 0;
      delete_midKey_293 <= 0;
      delete_success_294 <= 0;
      delete_test_295 <= 0;
      delete_next_296 <= 0;
      delete_root_297 <= 0;
      delete_isFree_298 <= 0;
      delete_next_299 <= 0;
      delete_root_300 <= 0;
      delete_isFree_301 <= 0;
      delete_index_302 <= 0;
      delete_size_303 <= 0;
      delete_isLeaf_304 <= 0;
      delete_nextFree_305 <= 0;
      delete_Key_0_306 <= 0;
      delete_KeyCompares_0_307 <= 0;
      delete_KeyCollapse_0_308 <= 0;
      delete_Data_0_309 <= 0;
      delete_Key_1_310 <= 0;
      delete_KeyCompares_1_311 <= 0;
      delete_KeyCollapse_1_312 <= 0;
      delete_Data_1_313 <= 0;
      delete_Key_2_314 <= 0;
      delete_KeyCompares_2_315 <= 0;
      delete_KeyCollapse_2_316 <= 0;
      delete_Data_2_317 <= 0;
      delete_Key_3_318 <= 0;
      delete_KeyCompares_3_319 <= 0;
      delete_KeyCollapse_3_320 <= 0;
      delete_Data_3_321 <= 0;
      delete_Found_322 <= 0;
      delete_Key_323 <= 0;
      delete_FoundKey_324 <= 0;
      delete_Data_325 <= 0;
      delete_BtreeIndex_326 <= 0;
      delete_StuckIndex_327 <= 0;
      delete_MergeSuccess_328 <= 0;
      delete_index_329 <= 0;
      delete_size_330 <= 0;
      delete_isLeaf_331 <= 0;
      delete_nextFree_332 <= 0;
      delete_Key_0_333 <= 0;
      delete_KeyCompares_0_334 <= 0;
      delete_KeyCollapse_0_335 <= 0;
      delete_Data_0_336 <= 0;
      delete_Key_1_337 <= 0;
      delete_KeyCompares_1_338 <= 0;
      delete_KeyCollapse_1_339 <= 0;
      delete_Data_1_340 <= 0;
      delete_Key_2_341 <= 0;
      delete_KeyCompares_2_342 <= 0;
      delete_KeyCollapse_2_343 <= 0;
      delete_Data_2_344 <= 0;
      delete_Key_3_345 <= 0;
      delete_KeyCompares_3_346 <= 0;
      delete_KeyCollapse_3_347 <= 0;
      delete_Data_3_348 <= 0;
      delete_Found_349 <= 0;
      delete_Key_350 <= 0;
      delete_FoundKey_351 <= 0;
      delete_Data_352 <= 0;
      delete_BtreeIndex_353 <= 0;
      delete_StuckIndex_354 <= 0;
      delete_MergeSuccess_355 <= 0;
      delete_childKey_356 <= 0;
      delete_size_357 <= 0;
      delete_childData_358 <= 0;
      delete_indexLeft_359 <= 0;
      delete_indexRight_360 <= 0;
      delete_midKey_361 <= 0;
      delete_success_362 <= 0;
      delete_test_363 <= 0;
      delete_next_364 <= 0;
      delete_root_365 <= 0;
      delete_isFree_366 <= 0;
      delete_index_367 <= 0;
      delete_size_368 <= 0;
      delete_isLeaf_369 <= 0;
      delete_nextFree_370 <= 0;
      delete_Key_0_371 <= 0;
      delete_KeyCompares_0_372 <= 0;
      delete_KeyCollapse_0_373 <= 0;
      delete_Data_0_374 <= 0;
      delete_Key_1_375 <= 0;
      delete_KeyCompares_1_376 <= 0;
      delete_KeyCollapse_1_377 <= 0;
      delete_Data_1_378 <= 0;
      delete_Key_2_379 <= 0;
      delete_KeyCompares_2_380 <= 0;
      delete_KeyCollapse_2_381 <= 0;
      delete_Data_2_382 <= 0;
      delete_Key_3_383 <= 0;
      delete_KeyCompares_3_384 <= 0;
      delete_KeyCollapse_3_385 <= 0;
      delete_Data_3_386 <= 0;
      delete_Found_387 <= 0;
      delete_Key_388 <= 0;
      delete_FoundKey_389 <= 0;
      delete_Data_390 <= 0;
      delete_BtreeIndex_391 <= 0;
      delete_StuckIndex_392 <= 0;
      delete_MergeSuccess_393 <= 0;
      delete_index_394 <= 0;
      delete_size_395 <= 0;
      delete_isLeaf_396 <= 0;
      delete_nextFree_397 <= 0;
      delete_Key_0_398 <= 0;
      delete_KeyCompares_0_399 <= 0;
      delete_KeyCollapse_0_400 <= 0;
      delete_Data_0_401 <= 0;
      delete_Key_1_402 <= 0;
      delete_KeyCompares_1_403 <= 0;
      delete_KeyCollapse_1_404 <= 0;
      delete_Data_1_405 <= 0;
      delete_Key_2_406 <= 0;
      delete_KeyCompares_2_407 <= 0;
      delete_KeyCollapse_2_408 <= 0;
      delete_Data_2_409 <= 0;
      delete_Key_3_410 <= 0;
      delete_KeyCompares_3_411 <= 0;
      delete_KeyCollapse_3_412 <= 0;
      delete_Data_3_413 <= 0;
      delete_Found_414 <= 0;
      delete_Key_415 <= 0;
      delete_FoundKey_416 <= 0;
      delete_Data_417 <= 0;
      delete_BtreeIndex_418 <= 0;
      delete_StuckIndex_419 <= 0;
      delete_MergeSuccess_420 <= 0;
      delete_childKey_421 <= 0;
      delete_size_422 <= 0;
      delete_childData_423 <= 0;
      delete_indexLeft_424 <= 0;
      delete_indexRight_425 <= 0;
      delete_midKey_426 <= 0;
      delete_success_427 <= 0;
      delete_test_428 <= 0;
      delete_next_429 <= 0;
      delete_root_430 <= 0;
      delete_isFree_431 <= 0;
      delete_index_432 <= 0;
      delete_size_433 <= 0;
      delete_isLeaf_434 <= 0;
      delete_nextFree_435 <= 0;
      delete_Key_0_436 <= 0;
      delete_KeyCompares_0_437 <= 0;
      delete_KeyCollapse_0_438 <= 0;
      delete_Data_0_439 <= 0;
      delete_Key_1_440 <= 0;
      delete_KeyCompares_1_441 <= 0;
      delete_KeyCollapse_1_442 <= 0;
      delete_Data_1_443 <= 0;
      delete_Key_2_444 <= 0;
      delete_KeyCompares_2_445 <= 0;
      delete_KeyCollapse_2_446 <= 0;
      delete_Data_2_447 <= 0;
      delete_Key_3_448 <= 0;
      delete_KeyCompares_3_449 <= 0;
      delete_KeyCollapse_3_450 <= 0;
      delete_Data_3_451 <= 0;
      delete_Found_452 <= 0;
      delete_Key_453 <= 0;
      delete_FoundKey_454 <= 0;
      delete_Data_455 <= 0;
      delete_BtreeIndex_456 <= 0;
      delete_StuckIndex_457 <= 0;
      delete_MergeSuccess_458 <= 0;
      delete_index_459 <= 0;
      delete_size_460 <= 0;
      delete_isLeaf_461 <= 0;
      delete_nextFree_462 <= 0;
      delete_Key_0_463 <= 0;
      delete_KeyCompares_0_464 <= 0;
      delete_KeyCollapse_0_465 <= 0;
      delete_Data_0_466 <= 0;
      delete_Key_1_467 <= 0;
      delete_KeyCompares_1_468 <= 0;
      delete_KeyCollapse_1_469 <= 0;
      delete_Data_1_470 <= 0;
      delete_Key_2_471 <= 0;
      delete_KeyCompares_2_472 <= 0;
      delete_KeyCollapse_2_473 <= 0;
      delete_Data_2_474 <= 0;
      delete_Key_3_475 <= 0;
      delete_KeyCompares_3_476 <= 0;
      delete_KeyCollapse_3_477 <= 0;
      delete_Data_3_478 <= 0;
      delete_Found_479 <= 0;
      delete_Key_480 <= 0;
      delete_FoundKey_481 <= 0;
      delete_Data_482 <= 0;
      delete_BtreeIndex_483 <= 0;
      delete_StuckIndex_484 <= 0;
      delete_MergeSuccess_485 <= 0;
      delete_childKey_486 <= 0;
      delete_childData_487 <= 0;
      delete_indexLeft_488 <= 0;
      delete_indexRight_489 <= 0;
      delete_midKey_490 <= 0;
      delete_success_491 <= 0;
      delete_test_492 <= 0;
      delete_next_493 <= 0;
      delete_root_494 <= 0;
      delete_isFree_495 <= 0;
      delete_index_496 <= 0;
      delete_size_497 <= 0;
      delete_isLeaf_498 <= 0;
      delete_nextFree_499 <= 0;
      delete_Key_0_500 <= 0;
      delete_KeyCompares_0_501 <= 0;
      delete_KeyCollapse_0_502 <= 0;
      delete_Data_0_503 <= 0;
      delete_Key_1_504 <= 0;
      delete_KeyCompares_1_505 <= 0;
      delete_KeyCollapse_1_506 <= 0;
      delete_Data_1_507 <= 0;
      delete_Key_2_508 <= 0;
      delete_KeyCompares_2_509 <= 0;
      delete_KeyCollapse_2_510 <= 0;
      delete_Data_2_511 <= 0;
      delete_Key_3_512 <= 0;
      delete_KeyCompares_3_513 <= 0;
      delete_KeyCollapse_3_514 <= 0;
      delete_Data_3_515 <= 0;
      delete_Found_516 <= 0;
      delete_Key_517 <= 0;
      delete_FoundKey_518 <= 0;
      delete_Data_519 <= 0;
      delete_BtreeIndex_520 <= 0;
      delete_StuckIndex_521 <= 0;
      delete_MergeSuccess_522 <= 0;
      delete_index_523 <= 0;
      delete_size_524 <= 0;
      delete_isLeaf_525 <= 0;
      delete_nextFree_526 <= 0;
      delete_Key_0_527 <= 0;
      delete_KeyCompares_0_528 <= 0;
      delete_KeyCollapse_0_529 <= 0;
      delete_Data_0_530 <= 0;
      delete_Key_1_531 <= 0;
      delete_KeyCompares_1_532 <= 0;
      delete_KeyCollapse_1_533 <= 0;
      delete_Data_1_534 <= 0;
      delete_Key_2_535 <= 0;
      delete_KeyCompares_2_536 <= 0;
      delete_KeyCollapse_2_537 <= 0;
      delete_Data_2_538 <= 0;
      delete_Key_3_539 <= 0;
      delete_KeyCompares_3_540 <= 0;
      delete_KeyCollapse_3_541 <= 0;
      delete_Data_3_542 <= 0;
      delete_Found_543 <= 0;
      delete_Key_544 <= 0;
      delete_FoundKey_545 <= 0;
      delete_Data_546 <= 0;
      delete_BtreeIndex_547 <= 0;
      delete_StuckIndex_548 <= 0;
      delete_MergeSuccess_549 <= 0;
      delete_childKey_550 <= 0;
      delete_leftChild_551 <= 0;
      delete_rightChild_552 <= 0;
      delete_childData_553 <= 0;
      delete_indexLeft_554 <= 0;
      delete_indexRight_555 <= 0;
      delete_midKey_556 <= 0;
      delete_success_557 <= 0;
      delete_test_558 <= 0;
      delete_next_559 <= 0;
      delete_root_560 <= 0;
      delete_isFree_561 <= 0;
      delete_index_562 <= 0;
      delete_size_563 <= 0;
      delete_isLeaf_564 <= 0;
      delete_nextFree_565 <= 0;
      delete_Key_0_566 <= 0;
      delete_KeyCompares_0_567 <= 0;
      delete_KeyCollapse_0_568 <= 0;
      delete_Data_0_569 <= 0;
      delete_Key_1_570 <= 0;
      delete_KeyCompares_1_571 <= 0;
      delete_KeyCollapse_1_572 <= 0;
      delete_Data_1_573 <= 0;
      delete_Key_2_574 <= 0;
      delete_KeyCompares_2_575 <= 0;
      delete_KeyCollapse_2_576 <= 0;
      delete_Data_2_577 <= 0;
      delete_Key_3_578 <= 0;
      delete_KeyCompares_3_579 <= 0;
      delete_KeyCollapse_3_580 <= 0;
      delete_Data_3_581 <= 0;
      delete_Found_582 <= 0;
      delete_Key_583 <= 0;
      delete_FoundKey_584 <= 0;
      delete_Data_585 <= 0;
      delete_BtreeIndex_586 <= 0;
      delete_StuckIndex_587 <= 0;
      delete_MergeSuccess_588 <= 0;
      delete_index_589 <= 0;
      delete_size_590 <= 0;
      delete_isLeaf_591 <= 0;
      delete_nextFree_592 <= 0;
      delete_Key_0_593 <= 0;
      delete_KeyCompares_0_594 <= 0;
      delete_KeyCollapse_0_595 <= 0;
      delete_Data_0_596 <= 0;
      delete_Key_1_597 <= 0;
      delete_KeyCompares_1_598 <= 0;
      delete_KeyCollapse_1_599 <= 0;
      delete_Data_1_600 <= 0;
      delete_Key_2_601 <= 0;
      delete_KeyCompares_2_602 <= 0;
      delete_KeyCollapse_2_603 <= 0;
      delete_Data_2_604 <= 0;
      delete_Key_3_605 <= 0;
      delete_KeyCompares_3_606 <= 0;
      delete_KeyCollapse_3_607 <= 0;
      delete_Data_3_608 <= 0;
      delete_Found_609 <= 0;
      delete_Key_610 <= 0;
      delete_FoundKey_611 <= 0;
      delete_Data_612 <= 0;
      delete_BtreeIndex_613 <= 0;
      delete_StuckIndex_614 <= 0;
      delete_MergeSuccess_615 <= 0;
      delete_childKey_616 <= 0;
      delete_childData_617 <= 0;
      delete_indexLeft_618 <= 0;
      delete_indexRight_619 <= 0;
      delete_midKey_620 <= 0;
      delete_success_621 <= 0;
      delete_test_622 <= 0;
      delete_next_623 <= 0;
      delete_root_624 <= 0;
      delete_isFree_625 <= 0;
      delete_index_626 <= 0;
      delete_size_627 <= 0;
      delete_isLeaf_628 <= 0;
      delete_nextFree_629 <= 0;
      delete_Key_0_630 <= 0;
      delete_KeyCompares_0_631 <= 0;
      delete_KeyCollapse_0_632 <= 0;
      delete_Data_0_633 <= 0;
      delete_Key_1_634 <= 0;
      delete_KeyCompares_1_635 <= 0;
      delete_KeyCollapse_1_636 <= 0;
      delete_Data_1_637 <= 0;
      delete_Key_2_638 <= 0;
      delete_KeyCompares_2_639 <= 0;
      delete_KeyCollapse_2_640 <= 0;
      delete_Data_2_641 <= 0;
      delete_Key_3_642 <= 0;
      delete_KeyCompares_3_643 <= 0;
      delete_KeyCollapse_3_644 <= 0;
      delete_Data_3_645 <= 0;
      delete_Found_646 <= 0;
      delete_Key_647 <= 0;
      delete_FoundKey_648 <= 0;
      delete_Data_649 <= 0;
      delete_BtreeIndex_650 <= 0;
      delete_StuckIndex_651 <= 0;
      delete_MergeSuccess_652 <= 0;
      delete_index_653 <= 0;
      delete_size_654 <= 0;
      delete_isLeaf_655 <= 0;
      delete_nextFree_656 <= 0;
      delete_Key_0_657 <= 0;
      delete_KeyCompares_0_658 <= 0;
      delete_KeyCollapse_0_659 <= 0;
      delete_Data_0_660 <= 0;
      delete_Key_1_661 <= 0;
      delete_KeyCompares_1_662 <= 0;
      delete_KeyCollapse_1_663 <= 0;
      delete_Data_1_664 <= 0;
      delete_Key_2_665 <= 0;
      delete_KeyCompares_2_666 <= 0;
      delete_KeyCollapse_2_667 <= 0;
      delete_Data_2_668 <= 0;
      delete_Key_3_669 <= 0;
      delete_KeyCompares_3_670 <= 0;
      delete_KeyCollapse_3_671 <= 0;
      delete_Data_3_672 <= 0;
      delete_Found_673 <= 0;
      delete_Key_674 <= 0;
      delete_FoundKey_675 <= 0;
      delete_Data_676 <= 0;
      delete_BtreeIndex_677 <= 0;
      delete_StuckIndex_678 <= 0;
      delete_MergeSuccess_679 <= 0;
      delete_childKey_680 <= 0;
      delete_leftChild_681 <= 0;
      delete_rightChild_682 <= 0;
      delete_childData_683 <= 0;
      delete_indexLeft_684 <= 0;
      delete_indexRight_685 <= 0;
      delete_midKey_686 <= 0;
      delete_success_687 <= 0;
      delete_test_688 <= 0;
      delete_next_689 <= 0;
      delete_root_690 <= 0;
      delete_isFree_691 <= 0;
      delete_index_692 <= 0;
      delete_size_693 <= 0;
      delete_isLeaf_694 <= 0;
      delete_nextFree_695 <= 0;
      delete_Key_0_696 <= 0;
      delete_KeyCompares_0_697 <= 0;
      delete_KeyCollapse_0_698 <= 0;
      delete_Data_0_699 <= 0;
      delete_Key_1_700 <= 0;
      delete_KeyCompares_1_701 <= 0;
      delete_KeyCollapse_1_702 <= 0;
      delete_Data_1_703 <= 0;
      delete_Key_2_704 <= 0;
      delete_KeyCompares_2_705 <= 0;
      delete_KeyCollapse_2_706 <= 0;
      delete_Data_2_707 <= 0;
      delete_Key_3_708 <= 0;
      delete_KeyCompares_3_709 <= 0;
      delete_KeyCollapse_3_710 <= 0;
      delete_Data_3_711 <= 0;
      delete_Found_712 <= 0;
      delete_Key_713 <= 0;
      delete_FoundKey_714 <= 0;
      delete_Data_715 <= 0;
      delete_BtreeIndex_716 <= 0;
      delete_StuckIndex_717 <= 0;
      delete_MergeSuccess_718 <= 0;
      delete_index_719 <= 0;
      delete_size_720 <= 0;
      delete_isLeaf_721 <= 0;
      delete_nextFree_722 <= 0;
      delete_Key_0_723 <= 0;
      delete_KeyCompares_0_724 <= 0;
      delete_KeyCollapse_0_725 <= 0;
      delete_Data_0_726 <= 0;
      delete_Key_1_727 <= 0;
      delete_KeyCompares_1_728 <= 0;
      delete_KeyCollapse_1_729 <= 0;
      delete_Data_1_730 <= 0;
      delete_Key_2_731 <= 0;
      delete_KeyCompares_2_732 <= 0;
      delete_KeyCollapse_2_733 <= 0;
      delete_Data_2_734 <= 0;
      delete_Key_3_735 <= 0;
      delete_KeyCompares_3_736 <= 0;
      delete_KeyCollapse_3_737 <= 0;
      delete_Data_3_738 <= 0;
      delete_Found_739 <= 0;
      delete_Key_740 <= 0;
      delete_FoundKey_741 <= 0;
      delete_Data_742 <= 0;
      delete_BtreeIndex_743 <= 0;
      delete_StuckIndex_744 <= 0;
      delete_MergeSuccess_745 <= 0;
      delete_childKey_746 <= 0;
      delete_childData_747 <= 0;
      delete_indexLeft_748 <= 0;
      delete_indexRight_749 <= 0;
      delete_midKey_750 <= 0;
      delete_success_751 <= 0;
      delete_test_752 <= 0;
      delete_next_753 <= 0;
      delete_root_754 <= 0;
      delete_isFree_755 <= 0;
      delete_index_756 <= 0;
      delete_size_757 <= 0;
      delete_isLeaf_758 <= 0;
      delete_nextFree_759 <= 0;
      delete_Key_0_760 <= 0;
      delete_KeyCompares_0_761 <= 0;
      delete_KeyCollapse_0_762 <= 0;
      delete_Data_0_763 <= 0;
      delete_Key_1_764 <= 0;
      delete_KeyCompares_1_765 <= 0;
      delete_KeyCollapse_1_766 <= 0;
      delete_Data_1_767 <= 0;
      delete_Key_2_768 <= 0;
      delete_KeyCompares_2_769 <= 0;
      delete_KeyCollapse_2_770 <= 0;
      delete_Data_2_771 <= 0;
      delete_Key_3_772 <= 0;
      delete_KeyCompares_3_773 <= 0;
      delete_KeyCollapse_3_774 <= 0;
      delete_Data_3_775 <= 0;
      delete_Found_776 <= 0;
      delete_Key_777 <= 0;
      delete_FoundKey_778 <= 0;
      delete_Data_779 <= 0;
      delete_BtreeIndex_780 <= 0;
      delete_StuckIndex_781 <= 0;
      delete_MergeSuccess_782 <= 0;
      delete_index_783 <= 0;
      delete_size_784 <= 0;
      delete_isLeaf_785 <= 0;
      delete_nextFree_786 <= 0;
      delete_Key_0_787 <= 0;
      delete_KeyCompares_0_788 <= 0;
      delete_KeyCollapse_0_789 <= 0;
      delete_Data_0_790 <= 0;
      delete_Key_1_791 <= 0;
      delete_KeyCompares_1_792 <= 0;
      delete_KeyCollapse_1_793 <= 0;
      delete_Data_1_794 <= 0;
      delete_Key_2_795 <= 0;
      delete_KeyCompares_2_796 <= 0;
      delete_KeyCollapse_2_797 <= 0;
      delete_Data_2_798 <= 0;
      delete_Key_3_799 <= 0;
      delete_KeyCompares_3_800 <= 0;
      delete_KeyCollapse_3_801 <= 0;
      delete_Data_3_802 <= 0;
      delete_Found_803 <= 0;
      delete_Key_804 <= 0;
      delete_FoundKey_805 <= 0;
      delete_Data_806 <= 0;
      delete_BtreeIndex_807 <= 0;
      delete_StuckIndex_808 <= 0;
      delete_MergeSuccess_809 <= 0;
      delete_childKey_810 <= 0;
      delete_leftChild_811 <= 0;
      delete_rightChild_812 <= 0;
      delete_childData_813 <= 0;
      delete_indexLeft_814 <= 0;
      delete_indexRight_815 <= 0;
      delete_midKey_816 <= 0;
      delete_success_817 <= 0;
      delete_test_818 <= 0;
      delete_next_819 <= 0;
      delete_root_820 <= 0;
      delete_isFree_821 <= 0;
      delete_index_822 <= 0;
      delete_size_823 <= 0;
      delete_isLeaf_824 <= 0;
      delete_nextFree_825 <= 0;
      delete_Key_0_826 <= 0;
      delete_KeyCompares_0_827 <= 0;
      delete_KeyCollapse_0_828 <= 0;
      delete_Data_0_829 <= 0;
      delete_Key_1_830 <= 0;
      delete_KeyCompares_1_831 <= 0;
      delete_KeyCollapse_1_832 <= 0;
      delete_Data_1_833 <= 0;
      delete_Key_2_834 <= 0;
      delete_KeyCompares_2_835 <= 0;
      delete_KeyCollapse_2_836 <= 0;
      delete_Data_2_837 <= 0;
      delete_Key_3_838 <= 0;
      delete_KeyCompares_3_839 <= 0;
      delete_KeyCollapse_3_840 <= 0;
      delete_Data_3_841 <= 0;
      delete_Found_842 <= 0;
      delete_Key_843 <= 0;
      delete_FoundKey_844 <= 0;
      delete_Data_845 <= 0;
      delete_BtreeIndex_846 <= 0;
      delete_StuckIndex_847 <= 0;
      delete_MergeSuccess_848 <= 0;
      delete_index_849 <= 0;
      delete_size_850 <= 0;
      delete_isLeaf_851 <= 0;
      delete_nextFree_852 <= 0;
      delete_Key_0_853 <= 0;
      delete_KeyCompares_0_854 <= 0;
      delete_KeyCollapse_0_855 <= 0;
      delete_Data_0_856 <= 0;
      delete_Key_1_857 <= 0;
      delete_KeyCompares_1_858 <= 0;
      delete_KeyCollapse_1_859 <= 0;
      delete_Data_1_860 <= 0;
      delete_Key_2_861 <= 0;
      delete_KeyCompares_2_862 <= 0;
      delete_KeyCollapse_2_863 <= 0;
      delete_Data_2_864 <= 0;
      delete_Key_3_865 <= 0;
      delete_KeyCompares_3_866 <= 0;
      delete_KeyCollapse_3_867 <= 0;
      delete_Data_3_868 <= 0;
      delete_Found_869 <= 0;
      delete_Key_870 <= 0;
      delete_FoundKey_871 <= 0;
      delete_Data_872 <= 0;
      delete_BtreeIndex_873 <= 0;
      delete_StuckIndex_874 <= 0;
      delete_MergeSuccess_875 <= 0;
      delete_childKey_876 <= 0;
      delete_childData_877 <= 0;
      delete_indexLeft_878 <= 0;
      delete_indexRight_879 <= 0;
      delete_midKey_880 <= 0;
      delete_success_881 <= 0;
      delete_test_882 <= 0;
      delete_next_883 <= 0;
      delete_root_884 <= 0;
      delete_isFree_885 <= 0;
      delete_index_886 <= 0;
      delete_size_887 <= 0;
      delete_isLeaf_888 <= 0;
      delete_nextFree_889 <= 0;
      delete_Key_0_890 <= 0;
      delete_KeyCompares_0_891 <= 0;
      delete_KeyCollapse_0_892 <= 0;
      delete_Data_0_893 <= 0;
      delete_Key_1_894 <= 0;
      delete_KeyCompares_1_895 <= 0;
      delete_KeyCollapse_1_896 <= 0;
      delete_Data_1_897 <= 0;
      delete_Key_2_898 <= 0;
      delete_KeyCompares_2_899 <= 0;
      delete_KeyCollapse_2_900 <= 0;
      delete_Data_2_901 <= 0;
      delete_Key_3_902 <= 0;
      delete_KeyCompares_3_903 <= 0;
      delete_KeyCollapse_3_904 <= 0;
      delete_Data_3_905 <= 0;
      delete_Found_906 <= 0;
      delete_Key_907 <= 0;
      delete_FoundKey_908 <= 0;
      delete_Data_909 <= 0;
      delete_BtreeIndex_910 <= 0;
      delete_StuckIndex_911 <= 0;
      delete_MergeSuccess_912 <= 0;
      delete_index_913 <= 0;
      delete_size_914 <= 0;
      delete_isLeaf_915 <= 0;
      delete_nextFree_916 <= 0;
      delete_Key_0_917 <= 0;
      delete_KeyCompares_0_918 <= 0;
      delete_KeyCollapse_0_919 <= 0;
      delete_Data_0_920 <= 0;
      delete_Key_1_921 <= 0;
      delete_KeyCompares_1_922 <= 0;
      delete_KeyCollapse_1_923 <= 0;
      delete_Data_1_924 <= 0;
      delete_Key_2_925 <= 0;
      delete_KeyCompares_2_926 <= 0;
      delete_KeyCollapse_2_927 <= 0;
      delete_Data_2_928 <= 0;
      delete_Key_3_929 <= 0;
      delete_KeyCompares_3_930 <= 0;
      delete_KeyCollapse_3_931 <= 0;
      delete_Data_3_932 <= 0;
      delete_Found_933 <= 0;
      delete_Key_934 <= 0;
      delete_FoundKey_935 <= 0;
      delete_Data_936 <= 0;
      delete_BtreeIndex_937 <= 0;
      delete_StuckIndex_938 <= 0;
      delete_MergeSuccess_939 <= 0;
      delete_childKey_940 <= 0;
      delete_leftChild_941 <= 0;
      delete_rightChild_942 <= 0;
      delete_childData_943 <= 0;
      delete_indexLeft_944 <= 0;
      delete_indexRight_945 <= 0;
      delete_midKey_946 <= 0;
      delete_success_947 <= 0;
      delete_test_948 <= 0;
      delete_next_949 <= 0;
      delete_root_950 <= 0;
      delete_isFree_951 <= 0;
      delete_index_952 <= 0;
      delete_size_953 <= 0;
      delete_isLeaf_954 <= 0;
      delete_nextFree_955 <= 0;
      delete_Key_0_956 <= 0;
      delete_KeyCompares_0_957 <= 0;
      delete_KeyCollapse_0_958 <= 0;
      delete_Data_0_959 <= 0;
      delete_Key_1_960 <= 0;
      delete_KeyCompares_1_961 <= 0;
      delete_KeyCollapse_1_962 <= 0;
      delete_Data_1_963 <= 0;
      delete_Key_2_964 <= 0;
      delete_KeyCompares_2_965 <= 0;
      delete_KeyCollapse_2_966 <= 0;
      delete_Data_2_967 <= 0;
      delete_Key_3_968 <= 0;
      delete_KeyCompares_3_969 <= 0;
      delete_KeyCollapse_3_970 <= 0;
      delete_Data_3_971 <= 0;
      delete_Found_972 <= 0;
      delete_Key_973 <= 0;
      delete_FoundKey_974 <= 0;
      delete_Data_975 <= 0;
      delete_BtreeIndex_976 <= 0;
      delete_StuckIndex_977 <= 0;
      delete_MergeSuccess_978 <= 0;
      delete_index_979 <= 0;
      delete_size_980 <= 0;
      delete_isLeaf_981 <= 0;
      delete_nextFree_982 <= 0;
      delete_Key_0_983 <= 0;
      delete_KeyCompares_0_984 <= 0;
      delete_KeyCollapse_0_985 <= 0;
      delete_Data_0_986 <= 0;
      delete_Key_1_987 <= 0;
      delete_KeyCompares_1_988 <= 0;
      delete_KeyCollapse_1_989 <= 0;
      delete_Data_1_990 <= 0;
      delete_Key_2_991 <= 0;
      delete_KeyCompares_2_992 <= 0;
      delete_KeyCollapse_2_993 <= 0;
      delete_Data_2_994 <= 0;
      delete_Key_3_995 <= 0;
      delete_KeyCompares_3_996 <= 0;
      delete_KeyCollapse_3_997 <= 0;
      delete_Data_3_998 <= 0;
      delete_Found_999 <= 0;
      delete_Key_1000 <= 0;
      delete_FoundKey_1001 <= 0;
      delete_Data_1002 <= 0;
      delete_BtreeIndex_1003 <= 0;
      delete_StuckIndex_1004 <= 0;
      delete_MergeSuccess_1005 <= 0;
      delete_childKey_1006 <= 0;
      delete_childData_1007 <= 0;
      delete_indexLeft_1008 <= 0;
      delete_indexRight_1009 <= 0;
      delete_midKey_1010 <= 0;
      delete_success_1011 <= 0;
      delete_test_1012 <= 0;
      delete_next_1013 <= 0;
      delete_root_1014 <= 0;
      delete_isFree_1015 <= 0;
      delete_index_1016 <= 0;
      delete_size_1017 <= 0;
      delete_isLeaf_1018 <= 0;
      delete_nextFree_1019 <= 0;
      delete_Key_0_1020 <= 0;
      delete_KeyCompares_0_1021 <= 0;
      delete_KeyCollapse_0_1022 <= 0;
      delete_Data_0_1023 <= 0;
      delete_Key_1_1024 <= 0;
      delete_KeyCompares_1_1025 <= 0;
      delete_KeyCollapse_1_1026 <= 0;
      delete_Data_1_1027 <= 0;
      delete_Key_2_1028 <= 0;
      delete_KeyCompares_2_1029 <= 0;
      delete_KeyCollapse_2_1030 <= 0;
      delete_Data_2_1031 <= 0;
      delete_Key_3_1032 <= 0;
      delete_KeyCompares_3_1033 <= 0;
      delete_KeyCollapse_3_1034 <= 0;
      delete_Data_3_1035 <= 0;
      delete_Found_1036 <= 0;
      delete_Key_1037 <= 0;
      delete_FoundKey_1038 <= 0;
      delete_Data_1039 <= 0;
      delete_BtreeIndex_1040 <= 0;
      delete_StuckIndex_1041 <= 0;
      delete_MergeSuccess_1042 <= 0;
      delete_index_1043 <= 0;
      delete_size_1044 <= 0;
      delete_isLeaf_1045 <= 0;
      delete_nextFree_1046 <= 0;
      delete_Key_0_1047 <= 0;
      delete_KeyCompares_0_1048 <= 0;
      delete_KeyCollapse_0_1049 <= 0;
      delete_Data_0_1050 <= 0;
      delete_Key_1_1051 <= 0;
      delete_KeyCompares_1_1052 <= 0;
      delete_KeyCollapse_1_1053 <= 0;
      delete_Data_1_1054 <= 0;
      delete_Key_2_1055 <= 0;
      delete_KeyCompares_2_1056 <= 0;
      delete_KeyCollapse_2_1057 <= 0;
      delete_Data_2_1058 <= 0;
      delete_Key_3_1059 <= 0;
      delete_KeyCompares_3_1060 <= 0;
      delete_KeyCollapse_3_1061 <= 0;
      delete_Data_3_1062 <= 0;
      delete_Found_1063 <= 0;
      delete_Key_1064 <= 0;
      delete_FoundKey_1065 <= 0;
      delete_Data_1066 <= 0;
      delete_BtreeIndex_1067 <= 0;
      delete_StuckIndex_1068 <= 0;
      delete_MergeSuccess_1069 <= 0;
      delete_childKey_1070 <= 0;
      delete_leftChild_1071 <= 0;
      delete_rightChild_1072 <= 0;
      delete_childData_1073 <= 0;
      delete_indexLeft_1074 <= 0;
      delete_indexRight_1075 <= 0;
      delete_midKey_1076 <= 0;
      delete_success_1077 <= 0;
      delete_test_1078 <= 0;
      delete_next_1079 <= 0;
      delete_root_1080 <= 0;
      delete_isFree_1081 <= 0;
      delete_index_1082 <= 0;
      delete_size_1083 <= 0;
      delete_isLeaf_1084 <= 0;
      delete_nextFree_1085 <= 0;
      delete_Key_0_1086 <= 0;
      delete_KeyCompares_0_1087 <= 0;
      delete_KeyCollapse_0_1088 <= 0;
      delete_Data_0_1089 <= 0;
      delete_Key_1_1090 <= 0;
      delete_KeyCompares_1_1091 <= 0;
      delete_KeyCollapse_1_1092 <= 0;
      delete_Data_1_1093 <= 0;
      delete_Key_2_1094 <= 0;
      delete_KeyCompares_2_1095 <= 0;
      delete_KeyCollapse_2_1096 <= 0;
      delete_Data_2_1097 <= 0;
      delete_Key_3_1098 <= 0;
      delete_KeyCompares_3_1099 <= 0;
      delete_KeyCollapse_3_1100 <= 0;
      delete_Data_3_1101 <= 0;
      delete_Found_1102 <= 0;
      delete_Key_1103 <= 0;
      delete_FoundKey_1104 <= 0;
      delete_Data_1105 <= 0;
      delete_BtreeIndex_1106 <= 0;
      delete_StuckIndex_1107 <= 0;
      delete_MergeSuccess_1108 <= 0;
      delete_index_1109 <= 0;
      delete_size_1110 <= 0;
      delete_isLeaf_1111 <= 0;
      delete_nextFree_1112 <= 0;
      delete_Key_0_1113 <= 0;
      delete_KeyCompares_0_1114 <= 0;
      delete_KeyCollapse_0_1115 <= 0;
      delete_Data_0_1116 <= 0;
      delete_Key_1_1117 <= 0;
      delete_KeyCompares_1_1118 <= 0;
      delete_KeyCollapse_1_1119 <= 0;
      delete_Data_1_1120 <= 0;
      delete_Key_2_1121 <= 0;
      delete_KeyCompares_2_1122 <= 0;
      delete_KeyCollapse_2_1123 <= 0;
      delete_Data_2_1124 <= 0;
      delete_Key_3_1125 <= 0;
      delete_KeyCompares_3_1126 <= 0;
      delete_KeyCollapse_3_1127 <= 0;
      delete_Data_3_1128 <= 0;
      delete_Found_1129 <= 0;
      delete_Key_1130 <= 0;
      delete_FoundKey_1131 <= 0;
      delete_Data_1132 <= 0;
      delete_BtreeIndex_1133 <= 0;
      delete_StuckIndex_1134 <= 0;
      delete_MergeSuccess_1135 <= 0;
      delete_childKey_1136 <= 0;
      delete_childData_1137 <= 0;
      delete_indexLeft_1138 <= 0;
      delete_indexRight_1139 <= 0;
      delete_midKey_1140 <= 0;
      delete_success_1141 <= 0;
      delete_test_1142 <= 0;
      delete_next_1143 <= 0;
      delete_root_1144 <= 0;
      delete_isFree_1145 <= 0;
      delete_index_1146 <= 0;
      delete_size_1147 <= 0;
      delete_isLeaf_1148 <= 0;
      delete_nextFree_1149 <= 0;
      delete_Key_0_1150 <= 0;
      delete_KeyCompares_0_1151 <= 0;
      delete_KeyCollapse_0_1152 <= 0;
      delete_Data_0_1153 <= 0;
      delete_Key_1_1154 <= 0;
      delete_KeyCompares_1_1155 <= 0;
      delete_KeyCollapse_1_1156 <= 0;
      delete_Data_1_1157 <= 0;
      delete_Key_2_1158 <= 0;
      delete_KeyCompares_2_1159 <= 0;
      delete_KeyCollapse_2_1160 <= 0;
      delete_Data_2_1161 <= 0;
      delete_Key_3_1162 <= 0;
      delete_KeyCompares_3_1163 <= 0;
      delete_KeyCollapse_3_1164 <= 0;
      delete_Data_3_1165 <= 0;
      delete_Found_1166 <= 0;
      delete_Key_1167 <= 0;
      delete_FoundKey_1168 <= 0;
      delete_Data_1169 <= 0;
      delete_BtreeIndex_1170 <= 0;
      delete_StuckIndex_1171 <= 0;
      delete_MergeSuccess_1172 <= 0;
      delete_index_1173 <= 0;
      delete_size_1174 <= 0;
      delete_isLeaf_1175 <= 0;
      delete_nextFree_1176 <= 0;
      delete_Key_0_1177 <= 0;
      delete_KeyCompares_0_1178 <= 0;
      delete_KeyCollapse_0_1179 <= 0;
      delete_Data_0_1180 <= 0;
      delete_Key_1_1181 <= 0;
      delete_KeyCompares_1_1182 <= 0;
      delete_KeyCollapse_1_1183 <= 0;
      delete_Data_1_1184 <= 0;
      delete_Key_2_1185 <= 0;
      delete_KeyCompares_2_1186 <= 0;
      delete_KeyCollapse_2_1187 <= 0;
      delete_Data_2_1188 <= 0;
      delete_Key_3_1189 <= 0;
      delete_KeyCompares_3_1190 <= 0;
      delete_KeyCollapse_3_1191 <= 0;
      delete_Data_3_1192 <= 0;
      delete_Found_1193 <= 0;
      delete_Key_1194 <= 0;
      delete_FoundKey_1195 <= 0;
      delete_Data_1196 <= 0;
      delete_BtreeIndex_1197 <= 0;
      delete_StuckIndex_1198 <= 0;
      delete_MergeSuccess_1199 <= 0;
      delete_childKey_1200 <= 0;
      delete_leftChild_1201 <= 0;
      delete_rightChild_1202 <= 0;
      delete_childData_1203 <= 0;
      delete_indexLeft_1204 <= 0;
      delete_indexRight_1205 <= 0;
      delete_midKey_1206 <= 0;
      delete_success_1207 <= 0;
      delete_test_1208 <= 0;
      delete_next_1209 <= 0;
      delete_root_1210 <= 0;
      delete_isFree_1211 <= 0;
      stuckIsLeaf_7_requestedAt <= -1;
      stuckIsLeaf_8_requestedAt <= -1;
      stuckIsFree_11_requestedAt <= -1;
      freeNext_9_requestedAt <= -1;
      freeNext_10_requestedAt <= -1;
      stuckSize_5_requestedAt <= -1;
      stuckSize_6_requestedAt <= -1;
      stuckKeys_1_requestedAt <= -1;
      stuckKeys_2_requestedAt <= -1;
      stuckData_3_requestedAt <= -1;
      stuckData_4_requestedAt <= -1;
    end
    else if (processCurrent == 6) begin
      case(delete_pc)
        0: begin
          delete_i_45 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0676:<init>|  Chip.java:0675:RegisterSet|  Btree.java:5306:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        1: begin
          case (delete_i_45)
            0: begin
              delete_k_46 <= 32;
              delete_i_45 <= delete_i_45+1;
            end
            1: begin
              delete_k_46 <= 31;
              delete_i_45 <= delete_i_45+1;
            end
            2: begin
              delete_k_46 <= 30;
              delete_i_45 <= delete_i_45+1;
            end
            3: begin
              delete_k_46 <= 29;
              delete_i_45 <= delete_i_45+1;
            end
            4: begin
              delete_k_46 <= 28;
              delete_i_45 <= delete_i_45+1;
            end
            5: begin
              delete_k_46 <= 27;
              delete_i_45 <= delete_i_45+1;
            end
            6: begin
              delete_k_46 <= 26;
              delete_i_45 <= delete_i_45+1;
            end
            7: begin
              delete_k_46 <= 25;
              delete_i_45 <= delete_i_45+1;
            end
            8: begin
              delete_k_46 <= 24;
              delete_i_45 <= delete_i_45+1;
            end
            9: begin
              delete_k_46 <= 23;
              delete_i_45 <= delete_i_45+1;
            end
            10: begin
              delete_k_46 <= 22;
              delete_i_45 <= delete_i_45+1;
            end
            11: begin
              delete_k_46 <= 21;
              delete_i_45 <= delete_i_45+1;
            end
            12: begin
              delete_k_46 <= 20;
              delete_i_45 <= delete_i_45+1;
            end
            13: begin
              delete_k_46 <= 19;
              delete_i_45 <= delete_i_45+1;
            end
            14: begin
              delete_k_46 <= 18;
              delete_i_45 <= delete_i_45+1;
            end
            15: begin
              delete_k_46 <= 17;
              delete_i_45 <= delete_i_45+1;
            end
            16: begin
              delete_k_46 <= 16;
              delete_i_45 <= delete_i_45+1;
            end
            17: begin
              delete_k_46 <= 15;
              delete_i_45 <= delete_i_45+1;
            end
            18: begin
              delete_k_46 <= 14;
              delete_i_45 <= delete_i_45+1;
            end
            19: begin
              delete_k_46 <= 13;
              delete_i_45 <= delete_i_45+1;
            end
            20: begin
              delete_k_46 <= 12;
              delete_i_45 <= delete_i_45+1;
            end
            21: begin
              delete_k_46 <= 11;
              delete_i_45 <= delete_i_45+1;
            end
            22: begin
              delete_k_46 <= 10;
              delete_i_45 <= delete_i_45+1;
            end
            23: begin
              delete_k_46 <= 9;
              delete_i_45 <= delete_i_45+1;
            end
            24: begin
              delete_k_46 <= 8;
              delete_i_45 <= delete_i_45+1;
            end
            25: begin
              delete_k_46 <= 7;
              delete_i_45 <= delete_i_45+1;
            end
            26: begin
              delete_k_46 <= 6;
              delete_i_45 <= delete_i_45+1;
            end
            27: begin
              delete_k_46 <= 5;
              delete_i_45 <= delete_i_45+1;
            end
            28: begin
              delete_k_46 <= 4;
              delete_i_45 <= delete_i_45+1;
            end
            29: begin
              delete_k_46 <= 3;
              delete_i_45 <= delete_i_45+1;
            end
            30: begin
              delete_k_46 <= 2;
              delete_i_45 <= delete_i_45+1;
            end
            31: begin
              delete_k_46 <= 1;
              delete_i_45 <= delete_i_45+1;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:5311:<init>|  Btree.java:5310:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        2: begin
          delete_BtreeIndex_72 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2250:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        3: begin
          delete_index_48 <= delete_BtreeIndex_72;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        4: begin
          delete_stuckSize_5_index_32 <= delete_index_48;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_48;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_48;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_48;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        5: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        6: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        7: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        8: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        9: begin
          delete_size_49 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_50 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_52 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_55 <= stuckData_stuckData_3_result_0;
          delete_Key_1_56 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_59 <= stuckData_stuckData_3_result_1;
          delete_Key_2_60 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_63 <= stuckData_stuckData_3_result_2;
          delete_Key_3_64 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_67 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        10: begin
          if (delete_isLeaf_50 == 0) begin
            delete_pc <= 17;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        11: begin
          delete_KeyCompares_0_53 <= delete_k_46 == delete_Key_0_52 && 0 < delete_size_49;
          delete_KeyCollapse_0_54 <= 0;
          delete_KeyCompares_1_57 <= delete_k_46 == delete_Key_1_56 && 1 < delete_size_49;
          delete_KeyCollapse_1_58 <= 1;
          delete_KeyCompares_2_61 <= delete_k_46 == delete_Key_2_60 && 2 < delete_size_49;
          delete_KeyCollapse_2_62 <= 2;
          delete_KeyCompares_3_65 <= delete_k_46 == delete_Key_3_64 && 3 < delete_size_49;
          delete_KeyCollapse_3_66 <= 3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0801:<init>|  Btree.java:0800:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        12: begin
          if (delete_KeyCompares_1_57) begin
            delete_KeyCompares_0_53 <= 1;
            delete_KeyCollapse_0_54 <= delete_KeyCollapse_1_58;
          end
          if (delete_KeyCompares_3_65) begin
            delete_KeyCompares_2_61 <= 1;
            delete_KeyCollapse_2_62 <= delete_KeyCollapse_3_66;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        13: begin
          if (delete_KeyCompares_2_61) begin
            delete_KeyCompares_0_53 <= 1;
            delete_KeyCollapse_0_54 <= delete_KeyCollapse_2_62;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        14: begin
          if (delete_KeyCompares_0_53) begin
            delete_Found_68 <= 1;
            case (delete_KeyCollapse_0_54)
              0: begin
                delete_StuckIndex_73 <= 0;
                delete_Key_69 <= delete_Key_0_52;
                delete_Data_71 <= delete_Data_0_55;
              end
              1: begin
                delete_StuckIndex_73 <= 1;
                delete_Key_69 <= delete_Key_1_56;
                delete_Data_71 <= delete_Data_1_59;
              end
              2: begin
                delete_StuckIndex_73 <= 2;
                delete_Key_69 <= delete_Key_2_60;
                delete_Data_71 <= delete_Data_2_63;
              end
              3: begin
                delete_StuckIndex_73 <= 3;
                delete_Key_69 <= delete_Key_3_64;
                delete_Data_71 <= delete_Data_3_67;
              end
            endcase
          end
          else begin
            delete_Found_68 <= 0;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0844:<init>|  Btree.java:0843:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        15: begin
          delete_pc <= 23;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2258:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        16: begin
          delete_pc <= 23;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        17: begin
          delete_KeyCompares_0_53 <= delete_k_46 <= delete_Key_0_52 && 0 < delete_size_49;
          delete_KeyCollapse_0_54 <= 0;
          delete_KeyCompares_1_57 <= delete_k_46 >  delete_Key_0_52 && delete_k_46 <= delete_Key_1_56 && 1 < delete_size_49;
          delete_KeyCollapse_1_58 <= 1;
          delete_KeyCompares_2_61 <= delete_k_46 >  delete_Key_1_56 && delete_k_46 <= delete_Key_2_60 && 2 < delete_size_49;
          delete_KeyCollapse_2_62 <= 2;
          delete_KeyCompares_3_65 <= delete_k_46 >  delete_Key_2_60 && delete_k_46 <= delete_Key_3_64 && 3 < delete_size_49;
          delete_KeyCollapse_3_66 <= 3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        18: begin
          if (delete_KeyCompares_1_57) begin
            delete_KeyCompares_0_53 <= 1;
            delete_KeyCollapse_0_54 <= delete_KeyCollapse_1_58;
          end
          if (delete_KeyCompares_3_65) begin
            delete_KeyCompares_2_61 <= 1;
            delete_KeyCollapse_2_62 <= delete_KeyCollapse_3_66;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        19: begin
          if (delete_KeyCompares_2_61) begin
            delete_KeyCompares_0_53 <= 1;
            delete_KeyCollapse_0_54 <= delete_KeyCollapse_2_62;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        20: begin
          if (delete_KeyCompares_0_53) begin
            delete_Found_68 <= 1;
            case (delete_KeyCollapse_0_54)
              0: begin
                delete_StuckIndex_73 <= 0;
                delete_FoundKey_70 <= delete_Key_0_52;
                delete_Data_71 <= delete_Data_0_55;
              end
              1: begin
                delete_StuckIndex_73 <= 1;
                delete_FoundKey_70 <= delete_Key_1_56;
                delete_Data_71 <= delete_Data_1_59;
              end
              2: begin
                delete_StuckIndex_73 <= 2;
                delete_FoundKey_70 <= delete_Key_2_60;
                delete_Data_71 <= delete_Data_2_63;
              end
              3: begin
                delete_StuckIndex_73 <= 3;
                delete_FoundKey_70 <= delete_Key_3_64;
                delete_Data_71 <= delete_Data_3_67;
              end
            endcase
          end
          else begin
            delete_Found_68 <= 0;
            case (delete_size_49)
              0: begin
                delete_StuckIndex_73 <= 0;
                delete_Data_71 <= delete_Data_0_55;
              end
              1: begin
                delete_StuckIndex_73 <= 1;
                delete_Data_71 <= delete_Data_1_59;
              end
              2: begin
                delete_StuckIndex_73 <= 2;
                delete_Data_71 <= delete_Data_2_63;
              end
              3: begin
                delete_StuckIndex_73 <= 3;
                delete_Data_71 <= delete_Data_3_67;
              end
            endcase
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        21: begin
          delete_BtreeIndex_72 <= delete_Data_71;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2262:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        22: begin
          delete_pc <= 3;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2263:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2622:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        23: begin
          if (delete_Found_68 == 0) begin
            delete_pc <= 853;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        24: begin
          delete_size_49 <= delete_size_49-1;
          case (delete_StuckIndex_73)
            0: begin
              delete_Key_69 <= delete_Key_0_52;
              delete_Data_71 <= delete_Data_0_55;
            end
            1: begin
              delete_Key_69 <= delete_Key_1_56;
              delete_Data_71 <= delete_Data_1_59;
            end
            2: begin
              delete_Key_69 <= delete_Key_2_60;
              delete_Data_71 <= delete_Data_2_63;
            end
            3: begin
              delete_Key_69 <= delete_Key_3_64;
              delete_Data_71 <= delete_Data_3_67;
            end
          endcase
          if (0>= delete_StuckIndex_73) begin
            delete_Key_0_52 <= delete_Key_1_56;
            delete_Data_0_55 <= delete_Data_1_59;
          end
          if (1>= delete_StuckIndex_73) begin
            delete_Key_1_56 <= delete_Key_2_60;
            delete_Data_1_59 <= delete_Data_2_63;
          end
          if (2>= delete_StuckIndex_73) begin
            delete_Key_2_60 <= delete_Key_3_64;
            delete_Data_2_63 <= delete_Data_3_67;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2626:<init>|  Btree.java:2625:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        25: begin
          delete_stuckSize_6_index_33 <= delete_index_48;
          delete_stuckSize_6_value_34 <= delete_size_49;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_48;
          delete_stuckKeys_2_value_22 <= delete_Key_0_52;
          delete_stuckKeys_2_value_23 <= delete_Key_1_56;
          delete_stuckKeys_2_value_24 <= delete_Key_2_60;
          delete_stuckKeys_2_value_25 <= delete_Key_3_64;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_48;
          delete_stuckData_4_value_28 <= delete_Data_0_55;
          delete_stuckData_4_value_29 <= delete_Data_1_59;
          delete_stuckData_4_value_30 <= delete_Data_2_63;
          delete_stuckData_4_value_31 <= delete_Data_3_67;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2633:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        26: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2633:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        27: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2633:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        28: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2633:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        29: begin
          delete_position_102 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2434:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        30: begin
          delete_index_75 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        31: begin
          delete_stuckSize_5_index_32 <= delete_index_75;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_75;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_75;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_75;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        32: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        33: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        34: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        35: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        36: begin
          delete_size_76 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_77 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_79 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_82 <= stuckData_stuckData_3_result_0;
          delete_Key_1_83 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_86 <= stuckData_stuckData_3_result_1;
          delete_Key_2_87 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_90 <= stuckData_stuckData_3_result_2;
          delete_Key_3_91 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_94 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        37: begin
          if (delete_isLeaf_77 == 0) begin
            delete_pc <= 40;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2439:<init>|  Btree.java:2438:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        38: begin
          delete_pc <= 852;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2440:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2439:<init>|  Btree.java:2438:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        39: begin
          delete_pc <= 40;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2439:<init>|  Btree.java:2438:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        40: begin
          delete_success_193 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1813:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        41: begin
          delete_index_107 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        42: begin
          delete_stuckSize_5_index_32 <= delete_index_107;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_107;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_107;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_107;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        43: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        44: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        45: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        46: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        47: begin
          delete_size_108 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_109 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_111 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_114 <= stuckData_stuckData_3_result_0;
          delete_Key_1_115 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_118 <= stuckData_stuckData_3_result_1;
          delete_Key_2_119 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_122 <= stuckData_stuckData_3_result_2;
          delete_Key_3_123 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_126 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        48: begin
          delete_test_194 <= delete_size_108==1 ? 1 : 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0785:<init>|  Chip.java:0785:Eq|  Btree.java:1816:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        49: begin
          if (delete_test_194 == 0) begin
            delete_pc <= 101;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0585:<init>|  Chip.java:0584:GOZero|  Btree.java:1817:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        50: begin
          delete_indexLeft_190 <= delete_Data_0_114;
          delete_indexRight_191 <= delete_Data_1_118;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1820:<init>|  Btree.java:1819:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        51: begin
          delete_index_134 <= delete_indexLeft_190;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        52: begin
          delete_stuckSize_5_index_32 <= delete_index_134;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_134;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_134;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_134;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        53: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        54: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        55: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        56: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        57: begin
          delete_size_135 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_136 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_138 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_141 <= stuckData_stuckData_3_result_0;
          delete_Key_1_142 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_145 <= stuckData_stuckData_3_result_1;
          delete_Key_2_146 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_149 <= stuckData_stuckData_3_result_2;
          delete_Key_3_150 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_153 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        58: begin
          delete_index_161 <= delete_indexRight_191;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        59: begin
          delete_stuckSize_5_index_32 <= delete_index_161;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_161;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_161;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_161;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        60: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        61: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        62: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        63: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        64: begin
          delete_size_162 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_163 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_165 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_168 <= stuckData_stuckData_3_result_0;
          delete_Key_1_169 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_172 <= stuckData_stuckData_3_result_1;
          delete_Key_2_173 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_176 <= stuckData_stuckData_3_result_2;
          delete_Key_3_177 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_180 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        65: begin
          if (delete_isLeaf_136 == 0) begin
            delete_pc <= 101;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        66: begin
          if (delete_isLeaf_163 == 0) begin
            delete_pc <= 100;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        67: begin
          delete_MergeSuccess_133 <= 0;
          case (delete_size_135)
            0: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                3: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                4: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                3: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1251:<init>|  Btree.java:1250:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        68: begin
          if (delete_MergeSuccess_133 == 0) begin
            delete_pc <= 72;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        69: begin
          delete_MergeSuccess_133 <= 0;
          case (delete_size_108)
            0: begin
              case (delete_size_135)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_0_111 <= delete_Key_0_138;
                  delete_Data_0_114 <= delete_Data_0_141;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_Key_0_111 <= delete_Key_0_138;
                  delete_Data_0_114 <= delete_Data_0_141;
                  delete_Key_1_115 <= delete_Key_1_142;
                  delete_Data_1_118 <= delete_Data_1_145;
                  delete_size_108 <= delete_size_108 + 2;
                  delete_MergeSuccess_133 <= 1;
                end
                3: begin
                  delete_Key_0_111 <= delete_Key_0_138;
                  delete_Data_0_114 <= delete_Data_0_141;
                  delete_Key_1_115 <= delete_Key_1_142;
                  delete_Data_1_118 <= delete_Data_1_145;
                  delete_Key_2_119 <= delete_Key_2_146;
                  delete_Data_2_122 <= delete_Data_2_149;
                  delete_size_108 <= delete_size_108 + 3;
                  delete_MergeSuccess_133 <= 1;
                end
                4: begin
                  delete_Key_0_111 <= delete_Key_0_138;
                  delete_Data_0_114 <= delete_Data_0_141;
                  delete_Key_1_115 <= delete_Key_1_142;
                  delete_Data_1_118 <= delete_Data_1_145;
                  delete_Key_2_119 <= delete_Key_2_146;
                  delete_Data_2_122 <= delete_Data_2_149;
                  delete_Key_3_123 <= delete_Key_3_150;
                  delete_Data_3_126 <= delete_Data_3_153;
                  delete_size_108 <= delete_size_108 + 4;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_135)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_1_115 <= delete_Key_0_138;
                  delete_Data_1_118 <= delete_Data_0_141;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_Key_1_115 <= delete_Key_0_138;
                  delete_Data_1_118 <= delete_Data_0_141;
                  delete_Key_2_119 <= delete_Key_1_142;
                  delete_Data_2_122 <= delete_Data_1_145;
                  delete_size_108 <= delete_size_108 + 2;
                  delete_MergeSuccess_133 <= 1;
                end
                3: begin
                  delete_Key_1_115 <= delete_Key_0_138;
                  delete_Data_1_118 <= delete_Data_0_141;
                  delete_Key_2_119 <= delete_Key_1_142;
                  delete_Data_2_122 <= delete_Data_1_145;
                  delete_Key_3_123 <= delete_Key_2_146;
                  delete_Data_3_126 <= delete_Data_2_149;
                  delete_size_108 <= delete_size_108 + 3;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_135)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_2_119 <= delete_Key_0_138;
                  delete_Data_2_122 <= delete_Data_0_141;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_Key_2_119 <= delete_Key_0_138;
                  delete_Data_2_122 <= delete_Data_0_141;
                  delete_Key_3_123 <= delete_Key_1_142;
                  delete_Data_3_126 <= delete_Data_1_145;
                  delete_size_108 <= delete_size_108 + 2;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_135)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_3_123 <= delete_Key_0_138;
                  delete_Data_3_126 <= delete_Data_0_141;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_135)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1279:Then|  Chip.java:0610:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        70: begin
          delete_MergeSuccess_133 <= 0;
          case (delete_size_108)
            0: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_0_111 <= delete_Key_0_165;
                  delete_Data_0_114 <= delete_Data_0_168;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_Key_0_111 <= delete_Key_0_165;
                  delete_Data_0_114 <= delete_Data_0_168;
                  delete_Key_1_115 <= delete_Key_1_169;
                  delete_Data_1_118 <= delete_Data_1_172;
                  delete_size_108 <= delete_size_108 + 2;
                  delete_MergeSuccess_133 <= 1;
                end
                3: begin
                  delete_Key_0_111 <= delete_Key_0_165;
                  delete_Data_0_114 <= delete_Data_0_168;
                  delete_Key_1_115 <= delete_Key_1_169;
                  delete_Data_1_118 <= delete_Data_1_172;
                  delete_Key_2_119 <= delete_Key_2_173;
                  delete_Data_2_122 <= delete_Data_2_176;
                  delete_size_108 <= delete_size_108 + 3;
                  delete_MergeSuccess_133 <= 1;
                end
                4: begin
                  delete_Key_0_111 <= delete_Key_0_165;
                  delete_Data_0_114 <= delete_Data_0_168;
                  delete_Key_1_115 <= delete_Key_1_169;
                  delete_Data_1_118 <= delete_Data_1_172;
                  delete_Key_2_119 <= delete_Key_2_173;
                  delete_Data_2_122 <= delete_Data_2_176;
                  delete_Key_3_123 <= delete_Key_3_177;
                  delete_Data_3_126 <= delete_Data_3_180;
                  delete_size_108 <= delete_size_108 + 4;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_1_115 <= delete_Key_0_165;
                  delete_Data_1_118 <= delete_Data_0_168;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_Key_1_115 <= delete_Key_0_165;
                  delete_Data_1_118 <= delete_Data_0_168;
                  delete_Key_2_119 <= delete_Key_1_169;
                  delete_Data_2_122 <= delete_Data_1_172;
                  delete_size_108 <= delete_size_108 + 2;
                  delete_MergeSuccess_133 <= 1;
                end
                3: begin
                  delete_Key_1_115 <= delete_Key_0_165;
                  delete_Data_1_118 <= delete_Data_0_168;
                  delete_Key_2_119 <= delete_Key_1_169;
                  delete_Data_2_122 <= delete_Data_1_172;
                  delete_Key_3_123 <= delete_Key_2_173;
                  delete_Data_3_126 <= delete_Data_2_176;
                  delete_size_108 <= delete_size_108 + 3;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_2_119 <= delete_Key_0_165;
                  delete_Data_2_122 <= delete_Data_0_168;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
                2: begin
                  delete_Key_2_119 <= delete_Key_0_165;
                  delete_Data_2_122 <= delete_Data_0_168;
                  delete_Key_3_123 <= delete_Key_1_169;
                  delete_Data_3_126 <= delete_Data_1_172;
                  delete_size_108 <= delete_size_108 + 2;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
                1: begin
                  delete_Key_3_123 <= delete_Key_0_165;
                  delete_Data_3_126 <= delete_Data_0_168;
                  delete_size_108 <= delete_size_108 + 1;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_162)
                0: begin
                  delete_size_108 <= delete_size_108 + 0;
                  delete_MergeSuccess_133 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1280:Then|  Chip.java:0610:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        71: begin
          delete_pc <= 72;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        72: begin
          if (delete_MergeSuccess_133 == 0) begin
            delete_pc <= 99;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        73: begin
          delete_isLeaf_109 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1840:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        74: begin
          delete_stuckSize_6_index_33 <= delete_index_107;
          delete_stuckSize_6_value_34 <= delete_size_108;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckIsLeaf_8_index_36 <= delete_index_107;
          delete_stuckIsLeaf_8_value_37 <= delete_isLeaf_109;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_107;
          delete_stuckKeys_2_value_22 <= delete_Key_0_111;
          delete_stuckKeys_2_value_23 <= delete_Key_1_115;
          delete_stuckKeys_2_value_24 <= delete_Key_2_119;
          delete_stuckKeys_2_value_25 <= delete_Key_3_123;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_107;
          delete_stuckData_4_value_28 <= delete_Data_0_114;
          delete_stuckData_4_value_29 <= delete_Data_1_118;
          delete_stuckData_4_value_30 <= delete_Data_2_122;
          delete_stuckData_4_value_31 <= delete_Data_3_126;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        75: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        76: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        77: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        78: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        79: begin
          delete_root_201 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        80: begin
          delete_freeNext_9_index_196 <= delete_root_201;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        81: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        82: begin
          delete_next_195 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_201;
          delete_freeNext_10_value_198 <= delete_indexLeft_190;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_202 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        83: begin
          delete_stuckIsFree_11_index_199 <= delete_indexLeft_190;
          delete_stuckIsFree_11_value_200 <= delete_isFree_202;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        84: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        85: begin
          delete_freeNext_10_index_197 <= delete_indexLeft_190;
          delete_freeNext_10_value_198 <= delete_next_195;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        86: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        87: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        88: begin
          delete_root_204 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        89: begin
          delete_freeNext_9_index_196 <= delete_root_204;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        90: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        91: begin
          delete_next_203 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_204;
          delete_freeNext_10_value_198 <= delete_indexRight_191;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_205 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        92: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_191;
          delete_stuckIsFree_11_value_200 <= delete_isFree_205;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        93: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        94: begin
          delete_freeNext_10_index_197 <= delete_indexRight_191;
          delete_freeNext_10_value_198 <= delete_next_203;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        95: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        96: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        97: begin
          delete_success_193 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1843:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        98: begin
          delete_pc <= 99;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        99: begin
          delete_pc <= 100;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        100: begin
          delete_pc <= 101;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        101: begin
          if (delete_success_193 == 0) begin
            delete_pc <= 104;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2444:<init>|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        102: begin
          delete_pc <= 852;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2445:Then|  Chip.java:0610:<init>|  Btree.java:2444:<init>|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        103: begin
          delete_pc <= 104;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2444:<init>|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        104: begin
          delete_index_206 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        105: begin
          delete_stuckSize_5_index_32 <= delete_index_206;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_206;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_206;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_206;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        106: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        107: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        108: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        109: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        110: begin
          delete_size_207 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_208 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_210 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_213 <= stuckData_stuckData_3_result_0;
          delete_Key_1_214 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_217 <= stuckData_stuckData_3_result_1;
          delete_Key_2_218 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_221 <= stuckData_stuckData_3_result_2;
          delete_Key_3_222 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_225 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        111: begin
          delete_success_294 <= 0;
          if (delete_size_207 != 1) begin
            delete_pc <= 157;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:2023:<init>|  Btree.java:2022:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        112: begin
          delete_midKey_293 <= delete_Key_0_210;
          delete_indexLeft_291 <= delete_Data_0_213;
          delete_indexRight_292 <= delete_Data_1_217;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2041:<init>|  Btree.java:2040:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        113: begin
          if (delete_isLeaf_235 == 0) begin
            delete_pc <= 115;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        114: begin
          delete_pc <= 157;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        115: begin
          if (delete_isLeaf_262 == 0) begin
            delete_pc <= 117;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        116: begin
          delete_pc <= 157;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        117: begin
          delete_index_233 <= delete_indexLeft_291;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        118: begin
          delete_stuckSize_5_index_32 <= delete_index_233;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_233;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_233;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_233;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        119: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        120: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        121: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        122: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        123: begin
          delete_size_234 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_235 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_237 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_240 <= stuckData_stuckData_3_result_0;
          delete_Key_1_241 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_244 <= stuckData_stuckData_3_result_1;
          delete_Key_2_245 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_248 <= stuckData_stuckData_3_result_2;
          delete_Key_3_249 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_252 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        124: begin
          delete_index_260 <= delete_indexRight_292;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        125: begin
          delete_stuckSize_5_index_32 <= delete_index_260;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_260;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_260;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_260;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        126: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        127: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        128: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        129: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        130: begin
          delete_size_261 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_262 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_264 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_267 <= stuckData_stuckData_3_result_0;
          delete_Key_1_268 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_271 <= stuckData_stuckData_3_result_1;
          delete_Key_2_272 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_275 <= stuckData_stuckData_3_result_2;
          delete_Key_3_276 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_279 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        131: begin
          delete_MergeSuccess_232 <= 0;
          case (delete_size_234)
            0: begin
              case (delete_size_261)
                0: begin
                  delete_Key_0_210 <= delete_midKey_293;
                  delete_Data_0_213 <= delete_Data_0_240;
                  delete_Data_1_217 <= delete_Data_0_267;
                  delete_size_207 <= 1;
                  delete_MergeSuccess_232 <= 1;
                end
                1: begin
                  delete_Key_0_210 <= delete_midKey_293;
                  delete_Data_0_213 <= delete_Data_0_240;
                  delete_Key_1_214 <= delete_Key_0_264;
                  delete_Data_1_217 <= delete_Data_0_267;
                  delete_Data_2_221 <= delete_Data_1_271;
                  delete_size_207 <= 2;
                  delete_MergeSuccess_232 <= 1;
                end
                2: begin
                  delete_Key_0_210 <= delete_midKey_293;
                  delete_Data_0_213 <= delete_Data_0_240;
                  delete_Key_1_214 <= delete_Key_0_264;
                  delete_Data_1_217 <= delete_Data_0_267;
                  delete_Key_2_218 <= delete_Key_1_268;
                  delete_Data_2_221 <= delete_Data_1_271;
                  delete_Data_3_225 <= delete_Data_2_275;
                  delete_size_207 <= 3;
                  delete_MergeSuccess_232 <= 1;
                end
                3: begin
                end
              endcase
            end
            1: begin
              case (delete_size_261)
                0: begin
                  delete_Key_0_210 <= delete_Key_0_237;
                  delete_Data_0_213 <= delete_Data_0_240;
                  delete_Key_1_214 <= delete_midKey_293;
                  delete_Data_1_217 <= delete_Data_1_244;
                  delete_Data_2_221 <= delete_Data_0_267;
                  delete_size_207 <= 2;
                  delete_MergeSuccess_232 <= 1;
                end
                1: begin
                  delete_Key_0_210 <= delete_Key_0_237;
                  delete_Data_0_213 <= delete_Data_0_240;
                  delete_Key_1_214 <= delete_midKey_293;
                  delete_Data_1_217 <= delete_Data_1_244;
                  delete_Key_2_218 <= delete_Key_0_264;
                  delete_Data_2_221 <= delete_Data_0_267;
                  delete_Data_3_225 <= delete_Data_1_271;
                  delete_size_207 <= 3;
                  delete_MergeSuccess_232 <= 1;
                end
                2: begin
                end
              endcase
            end
            2: begin
              case (delete_size_261)
                0: begin
                  delete_Key_0_210 <= delete_Key_0_237;
                  delete_Data_0_213 <= delete_Data_0_240;
                  delete_Key_1_214 <= delete_Key_1_241;
                  delete_Data_1_217 <= delete_Data_1_244;
                  delete_Key_2_218 <= delete_midKey_293;
                  delete_Data_2_221 <= delete_Data_2_248;
                  delete_Data_3_225 <= delete_Data_0_267;
                  delete_size_207 <= 3;
                  delete_MergeSuccess_232 <= 1;
                end
                1: begin
                end
              endcase
            end
            3: begin
              case (delete_size_261)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1329:<init>|  Btree.java:1328:mergeButOne|  Btree.java:2059:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        132: begin
          if (delete_MergeSuccess_232 == 0) begin
            delete_pc <= 157;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        133: begin
          delete_stuckSize_6_index_33 <= delete_index_206;
          delete_stuckSize_6_value_34 <= delete_size_207;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_206;
          delete_stuckKeys_2_value_22 <= delete_Key_0_210;
          delete_stuckKeys_2_value_23 <= delete_Key_1_214;
          delete_stuckKeys_2_value_24 <= delete_Key_2_218;
          delete_stuckKeys_2_value_25 <= delete_Key_3_222;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_206;
          delete_stuckData_4_value_28 <= delete_Data_0_213;
          delete_stuckData_4_value_29 <= delete_Data_1_217;
          delete_stuckData_4_value_30 <= delete_Data_2_221;
          delete_stuckData_4_value_31 <= delete_Data_3_225;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        134: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        135: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        136: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        137: begin
          delete_root_297 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        138: begin
          delete_freeNext_9_index_196 <= delete_root_297;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        139: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        140: begin
          delete_next_296 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_297;
          delete_freeNext_10_value_198 <= delete_indexLeft_291;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_298 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        141: begin
          delete_stuckIsFree_11_index_199 <= delete_indexLeft_291;
          delete_stuckIsFree_11_value_200 <= delete_isFree_298;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        142: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        143: begin
          delete_freeNext_10_index_197 <= delete_indexLeft_291;
          delete_freeNext_10_value_198 <= delete_next_296;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        144: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        145: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        146: begin
          delete_root_300 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        147: begin
          delete_freeNext_9_index_196 <= delete_root_300;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        148: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        149: begin
          delete_next_299 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_300;
          delete_freeNext_10_value_198 <= delete_indexRight_292;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_301 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        150: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_292;
          delete_stuckIsFree_11_value_200 <= delete_isFree_301;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        151: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        152: begin
          delete_freeNext_10_index_197 <= delete_indexRight_292;
          delete_freeNext_10_value_198 <= delete_next_299;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        153: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        154: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        155: begin
          delete_success_294 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2064:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        156: begin
          delete_pc <= 157;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        157: begin
          if (delete_success_294 == 0) begin
            delete_pc <= 166;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        158: begin
          delete_index_75 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        159: begin
          delete_stuckSize_5_index_32 <= delete_index_75;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_75;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_75;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_75;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        160: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        161: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        162: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        163: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        164: begin
          delete_size_76 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_77 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_79 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_82 <= stuckData_stuckData_3_result_0;
          delete_Key_1_83 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_86 <= stuckData_stuckData_3_result_1;
          delete_Key_2_87 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_90 <= stuckData_stuckData_3_result_2;
          delete_Key_3_91 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_94 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        165: begin
          delete_pc <= 166;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        166: begin
          delete_success_362 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1941:<init>|  Btree.java:1940:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        167: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 209;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1949:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        168: begin
          delete_size_357 <= delete_size_76;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1950:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        169: begin
          case (delete_size_357)
            1: begin
              delete_indexLeft_359 <= delete_Data_0_82;
              delete_indexRight_360 <= delete_Data_1_86;
            end
            2: begin
              delete_indexLeft_359 <= delete_Data_1_86;
              delete_indexRight_360 <= delete_Data_2_90;
            end
            3: begin
              delete_indexLeft_359 <= delete_Data_2_90;
              delete_indexRight_360 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1953:<init>|  Btree.java:1952:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        170: begin
          delete_index_302 <= delete_indexLeft_359;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        171: begin
          delete_stuckSize_5_index_32 <= delete_index_302;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_302;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_302;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_302;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        172: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        173: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        174: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        175: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        176: begin
          delete_size_303 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_304 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_306 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_309 <= stuckData_stuckData_3_result_0;
          delete_Key_1_310 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_313 <= stuckData_stuckData_3_result_1;
          delete_Key_2_314 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_317 <= stuckData_stuckData_3_result_2;
          delete_Key_3_318 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_321 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        177: begin
          delete_index_329 <= delete_indexRight_360;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        178: begin
          delete_stuckSize_5_index_32 <= delete_index_329;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_329;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_329;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_329;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        179: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        180: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        181: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        182: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        183: begin
          delete_size_330 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_331 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_333 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_336 <= stuckData_stuckData_3_result_0;
          delete_Key_1_337 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_340 <= stuckData_stuckData_3_result_1;
          delete_Key_2_341 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_344 <= stuckData_stuckData_3_result_2;
          delete_Key_3_345 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_348 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        184: begin
          if (delete_isLeaf_304 == 0) begin
            delete_pc <= 209;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        185: begin
          if (delete_isLeaf_331 == 0) begin
            delete_pc <= 208;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        186: begin
          delete_MergeSuccess_328 <= 0;
          case (delete_size_303)
            0: begin
              case (delete_size_330)
                0: begin
                  delete_size_303 <= delete_size_303 + 0;
                  delete_MergeSuccess_328 <= 1;
                end
                1: begin
                  delete_Key_0_306 <= delete_Key_0_333;
                  delete_Data_0_309 <= delete_Data_0_336;
                  delete_size_303 <= delete_size_303 + 1;
                  delete_MergeSuccess_328 <= 1;
                end
                2: begin
                  delete_Key_0_306 <= delete_Key_0_333;
                  delete_Data_0_309 <= delete_Data_0_336;
                  delete_Key_1_310 <= delete_Key_1_337;
                  delete_Data_1_313 <= delete_Data_1_340;
                  delete_size_303 <= delete_size_303 + 2;
                  delete_MergeSuccess_328 <= 1;
                end
                3: begin
                  delete_Key_0_306 <= delete_Key_0_333;
                  delete_Data_0_309 <= delete_Data_0_336;
                  delete_Key_1_310 <= delete_Key_1_337;
                  delete_Data_1_313 <= delete_Data_1_340;
                  delete_Key_2_314 <= delete_Key_2_341;
                  delete_Data_2_317 <= delete_Data_2_344;
                  delete_size_303 <= delete_size_303 + 3;
                  delete_MergeSuccess_328 <= 1;
                end
                4: begin
                  delete_Key_0_306 <= delete_Key_0_333;
                  delete_Data_0_309 <= delete_Data_0_336;
                  delete_Key_1_310 <= delete_Key_1_337;
                  delete_Data_1_313 <= delete_Data_1_340;
                  delete_Key_2_314 <= delete_Key_2_341;
                  delete_Data_2_317 <= delete_Data_2_344;
                  delete_Key_3_318 <= delete_Key_3_345;
                  delete_Data_3_321 <= delete_Data_3_348;
                  delete_size_303 <= delete_size_303 + 4;
                  delete_MergeSuccess_328 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_330)
                0: begin
                  delete_size_303 <= delete_size_303 + 0;
                  delete_MergeSuccess_328 <= 1;
                end
                1: begin
                  delete_Key_1_310 <= delete_Key_0_333;
                  delete_Data_1_313 <= delete_Data_0_336;
                  delete_size_303 <= delete_size_303 + 1;
                  delete_MergeSuccess_328 <= 1;
                end
                2: begin
                  delete_Key_1_310 <= delete_Key_0_333;
                  delete_Data_1_313 <= delete_Data_0_336;
                  delete_Key_2_314 <= delete_Key_1_337;
                  delete_Data_2_317 <= delete_Data_1_340;
                  delete_size_303 <= delete_size_303 + 2;
                  delete_MergeSuccess_328 <= 1;
                end
                3: begin
                  delete_Key_1_310 <= delete_Key_0_333;
                  delete_Data_1_313 <= delete_Data_0_336;
                  delete_Key_2_314 <= delete_Key_1_337;
                  delete_Data_2_317 <= delete_Data_1_340;
                  delete_Key_3_318 <= delete_Key_2_341;
                  delete_Data_3_321 <= delete_Data_2_344;
                  delete_size_303 <= delete_size_303 + 3;
                  delete_MergeSuccess_328 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_330)
                0: begin
                  delete_size_303 <= delete_size_303 + 0;
                  delete_MergeSuccess_328 <= 1;
                end
                1: begin
                  delete_Key_2_314 <= delete_Key_0_333;
                  delete_Data_2_317 <= delete_Data_0_336;
                  delete_size_303 <= delete_size_303 + 1;
                  delete_MergeSuccess_328 <= 1;
                end
                2: begin
                  delete_Key_2_314 <= delete_Key_0_333;
                  delete_Data_2_317 <= delete_Data_0_336;
                  delete_Key_3_318 <= delete_Key_1_337;
                  delete_Data_3_321 <= delete_Data_1_340;
                  delete_size_303 <= delete_size_303 + 2;
                  delete_MergeSuccess_328 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_330)
                0: begin
                  delete_size_303 <= delete_size_303 + 0;
                  delete_MergeSuccess_328 <= 1;
                end
                1: begin
                  delete_Key_3_318 <= delete_Key_0_333;
                  delete_Data_3_321 <= delete_Data_0_336;
                  delete_size_303 <= delete_size_303 + 1;
                  delete_MergeSuccess_328 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_330)
                0: begin
                  delete_size_303 <= delete_size_303 + 0;
                  delete_MergeSuccess_328 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1974:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        187: begin
          if (delete_MergeSuccess_328 == 0) begin
            delete_pc <= 207;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        188: begin
          delete_size_76 <= delete_size_76-1;
          delete_success_362 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1978:<init>|  Btree.java:1977:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        189: begin
          delete_stuckSize_6_index_33 <= delete_index_302;
          delete_stuckSize_6_value_34 <= delete_size_303;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_302;
          delete_stuckKeys_2_value_22 <= delete_Key_0_306;
          delete_stuckKeys_2_value_23 <= delete_Key_1_310;
          delete_stuckKeys_2_value_24 <= delete_Key_2_314;
          delete_stuckKeys_2_value_25 <= delete_Key_3_318;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_302;
          delete_stuckData_4_value_28 <= delete_Data_0_309;
          delete_stuckData_4_value_29 <= delete_Data_1_313;
          delete_stuckData_4_value_30 <= delete_Data_2_317;
          delete_stuckData_4_value_31 <= delete_Data_3_321;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        190: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        191: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        192: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        193: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        194: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        195: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        196: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        197: begin
          delete_root_365 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        198: begin
          delete_freeNext_9_index_196 <= delete_root_365;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        199: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        200: begin
          delete_next_364 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_365;
          delete_freeNext_10_value_198 <= delete_indexRight_360;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_366 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        201: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_360;
          delete_stuckIsFree_11_value_200 <= delete_isFree_366;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        202: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        203: begin
          delete_freeNext_10_index_197 <= delete_indexRight_360;
          delete_freeNext_10_value_198 <= delete_next_364;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        204: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        205: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        206: begin
          delete_pc <= 207;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        207: begin
          delete_pc <= 208;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        208: begin
          delete_pc <= 209;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        209: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 254;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2183:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        210: begin
          delete_success_427 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2184:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        211: begin
          delete_size_422 <= delete_size_76;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2185:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        212: begin
          case (delete_size_422)
            1: begin
              delete_indexLeft_424 <= delete_Data_0_82;
              delete_indexRight_425 <= delete_Data_1_86;
            end
            2: begin
              delete_indexLeft_424 <= delete_Data_1_86;
              delete_indexRight_425 <= delete_Data_2_90;
            end
            3: begin
              delete_indexLeft_424 <= delete_Data_2_90;
              delete_indexRight_425 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2188:<init>|  Btree.java:2187:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        213: begin
          delete_index_367 <= delete_indexLeft_424;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        214: begin
          delete_stuckSize_5_index_32 <= delete_index_367;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_367;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_367;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_367;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        215: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        216: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        217: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        218: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        219: begin
          delete_size_368 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_369 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_371 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_374 <= stuckData_stuckData_3_result_0;
          delete_Key_1_375 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_378 <= stuckData_stuckData_3_result_1;
          delete_Key_2_379 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_382 <= stuckData_stuckData_3_result_2;
          delete_Key_3_383 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_386 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        220: begin
          delete_index_394 <= delete_indexRight_425;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        221: begin
          delete_stuckSize_5_index_32 <= delete_index_394;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_394;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_394;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_394;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        222: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        223: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        224: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        225: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        226: begin
          delete_size_395 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_396 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_398 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_401 <= stuckData_stuckData_3_result_0;
          delete_Key_1_402 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_405 <= stuckData_stuckData_3_result_1;
          delete_Key_2_406 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_409 <= stuckData_stuckData_3_result_2;
          delete_Key_3_410 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_413 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        227: begin
          if (delete_isLeaf_369 == 0) begin
            delete_pc <= 229;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        228: begin
          delete_pc <= 254;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        229: begin
          if (delete_isLeaf_396 == 0) begin
            delete_pc <= 231;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        230: begin
          delete_pc <= 254;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        231: begin
          case (delete_size_76)
            1: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            2: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            3: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            4: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_size_76 <= delete_size_76-1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0452:<init>|  Btree.java:0451:Pop|  Btree.java:2209:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        232: begin
          delete_MergeSuccess_393 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2210:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        233: begin
          case (delete_size_368)
            0: begin
              case (delete_size_395)
                0: begin
                  delete_Key_0_371 <= delete_Key_96;
                  delete_Data_1_378 <= delete_Data_0_401;
                  delete_size_368 <= delete_size_368 + 1;
                  delete_MergeSuccess_393 <= 1;
                end
                1: begin
                  delete_Key_0_371 <= delete_Key_96;
                  delete_Key_1_375 <= delete_Key_0_398;
                  delete_Data_1_378 <= delete_Data_0_401;
                  delete_Data_2_382 <= delete_Data_1_405;
                  delete_size_368 <= delete_size_368 + 2;
                  delete_MergeSuccess_393 <= 1;
                end
                2: begin
                  delete_Key_0_371 <= delete_Key_96;
                  delete_Key_1_375 <= delete_Key_0_398;
                  delete_Data_1_378 <= delete_Data_0_401;
                  delete_Key_2_379 <= delete_Key_1_402;
                  delete_Data_2_382 <= delete_Data_1_405;
                  delete_Data_3_386 <= delete_Data_2_409;
                  delete_size_368 <= delete_size_368 + 3;
                  delete_MergeSuccess_393 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_395)
                0: begin
                  delete_Key_1_375 <= delete_Key_96;
                  delete_Data_2_382 <= delete_Data_0_401;
                  delete_size_368 <= delete_size_368 + 1;
                  delete_MergeSuccess_393 <= 1;
                end
                1: begin
                  delete_Key_1_375 <= delete_Key_96;
                  delete_Key_2_379 <= delete_Key_0_398;
                  delete_Data_2_382 <= delete_Data_0_401;
                  delete_Data_3_386 <= delete_Data_1_405;
                  delete_size_368 <= delete_size_368 + 2;
                  delete_MergeSuccess_393 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_395)
                0: begin
                  delete_Key_2_379 <= delete_Key_96;
                  delete_Data_3_386 <= delete_Data_0_401;
                  delete_size_368 <= delete_size_368 + 1;
                  delete_MergeSuccess_393 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_395)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_395)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2210:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        234: begin
          if (delete_MergeSuccess_393 == 0) begin
            delete_pc <= 254;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        235: begin
          delete_success_427 <= 1;
          case (delete_size_76)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_424;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_424;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_424;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_424;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2214:<init>|  Btree.java:2213:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        236: begin
          delete_stuckSize_6_index_33 <= delete_index_367;
          delete_stuckSize_6_value_34 <= delete_size_368;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_367;
          delete_stuckKeys_2_value_22 <= delete_Key_0_371;
          delete_stuckKeys_2_value_23 <= delete_Key_1_375;
          delete_stuckKeys_2_value_24 <= delete_Key_2_379;
          delete_stuckKeys_2_value_25 <= delete_Key_3_383;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_367;
          delete_stuckData_4_value_28 <= delete_Data_0_374;
          delete_stuckData_4_value_29 <= delete_Data_1_378;
          delete_stuckData_4_value_30 <= delete_Data_2_382;
          delete_stuckData_4_value_31 <= delete_Data_3_386;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        237: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        238: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        239: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        240: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        241: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        242: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        243: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        244: begin
          delete_root_430 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        245: begin
          delete_freeNext_9_index_196 <= delete_root_430;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        246: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        247: begin
          delete_next_429 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_430;
          delete_freeNext_10_value_198 <= delete_indexRight_425;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_431 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        248: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_425;
          delete_stuckIsFree_11_value_200 <= delete_isFree_431;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        249: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        250: begin
          delete_freeNext_10_index_197 <= delete_indexRight_425;
          delete_freeNext_10_value_198 <= delete_next_429;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        251: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        252: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        253: begin
          delete_pc <= 254;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        254: begin
          delete_index_75 <= delete_position_102;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        255: begin
          delete_stuckSize_5_index_32 <= delete_index_75;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_75;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_75;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_75;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        256: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        257: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        258: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        259: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        260: begin
          delete_size_76 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_77 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_79 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_82 <= stuckData_stuckData_3_result_0;
          delete_Key_1_83 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_86 <= stuckData_stuckData_3_result_1;
          delete_Key_2_87 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_90 <= stuckData_stuckData_3_result_2;
          delete_Key_3_91 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_94 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        261: begin
          delete_KeyCompares_0_80 <= delete_k_46 <= delete_Key_0_79 && 0 < delete_size_76;
          delete_KeyCollapse_0_81 <= 0;
          delete_KeyCompares_1_84 <= delete_k_46 >  delete_Key_0_79 && delete_k_46 <= delete_Key_1_83 && 1 < delete_size_76;
          delete_KeyCollapse_1_85 <= 1;
          delete_KeyCompares_2_88 <= delete_k_46 >  delete_Key_1_83 && delete_k_46 <= delete_Key_2_87 && 2 < delete_size_76;
          delete_KeyCollapse_2_89 <= 2;
          delete_KeyCompares_3_92 <= delete_k_46 >  delete_Key_2_87 && delete_k_46 <= delete_Key_3_91 && 3 < delete_size_76;
          delete_KeyCollapse_3_93 <= 3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2460:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        262: begin
          if (delete_KeyCompares_1_84) begin
            delete_KeyCompares_0_80 <= 1;
            delete_KeyCollapse_0_81 <= delete_KeyCollapse_1_85;
          end
          if (delete_KeyCompares_3_92) begin
            delete_KeyCompares_2_88 <= 1;
            delete_KeyCollapse_2_89 <= delete_KeyCollapse_3_93;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2460:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        263: begin
          if (delete_KeyCompares_2_88) begin
            delete_KeyCompares_0_80 <= 1;
            delete_KeyCollapse_0_81 <= delete_KeyCollapse_2_89;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2460:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        264: begin
          if (delete_KeyCompares_0_80) begin
            delete_Found_95 <= 1;
            case (delete_KeyCollapse_0_81)
              0: begin
                delete_StuckIndex_100 <= 0;
                delete_FoundKey_97 <= delete_Key_0_79;
                delete_Data_98 <= delete_Data_0_82;
              end
              1: begin
                delete_StuckIndex_100 <= 1;
                delete_FoundKey_97 <= delete_Key_1_83;
                delete_Data_98 <= delete_Data_1_86;
              end
              2: begin
                delete_StuckIndex_100 <= 2;
                delete_FoundKey_97 <= delete_Key_2_87;
                delete_Data_98 <= delete_Data_2_90;
              end
              3: begin
                delete_StuckIndex_100 <= 3;
                delete_FoundKey_97 <= delete_Key_3_91;
                delete_Data_98 <= delete_Data_3_94;
              end
            endcase
          end
          else begin
            delete_Found_95 <= 0;
            case (delete_size_76)
              0: begin
                delete_StuckIndex_100 <= 0;
                delete_Data_98 <= delete_Data_0_82;
              end
              1: begin
                delete_StuckIndex_100 <= 1;
                delete_Data_98 <= delete_Data_1_86;
              end
              2: begin
                delete_StuckIndex_100 <= 2;
                delete_Data_98 <= delete_Data_2_90;
              end
              3: begin
                delete_StuckIndex_100 <= 3;
                delete_Data_98 <= delete_Data_3_94;
              end
            endcase
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2460:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        265: begin
          if (delete_Found_95 == 0) begin
            delete_pc <= 731;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        266: begin
          if (delete_StuckIndex_100 == 0) begin
            delete_pc <= 548;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        267: begin
          delete_index1_104 <= delete_StuckIndex_100;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2466:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        268: begin
          delete_index1_104 <= delete_index1_104+1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0806:<init>|  Chip.java:0805:Inc|  Btree.java:2467:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        269: begin
          delete_within_105 <= delete_index1_104< delete_size_76 ? 1 : 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0781:<init>|  Chip.java:0781:Lt|  Btree.java:2469:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        270: begin
          if (delete_within_105 == 0) begin
            delete_pc <= 363;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        271: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 315;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        272: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_488 <= delete_Data_0_82;
              delete_indexRight_489 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_488 <= delete_Data_1_86;
              delete_indexRight_489 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_488 <= delete_Data_2_90;
              delete_indexRight_489 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        273: begin
          delete_index_432 <= delete_indexLeft_488;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        274: begin
          delete_stuckSize_5_index_32 <= delete_index_432;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_432;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_432;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_432;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        275: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        276: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        277: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        278: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        279: begin
          delete_size_433 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_434 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_436 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_439 <= stuckData_stuckData_3_result_0;
          delete_Key_1_440 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_443 <= stuckData_stuckData_3_result_1;
          delete_Key_2_444 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_447 <= stuckData_stuckData_3_result_2;
          delete_Key_3_448 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_451 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        280: begin
          delete_index_459 <= delete_indexRight_489;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        281: begin
          delete_stuckSize_5_index_32 <= delete_index_459;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_459;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_459;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_459;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        282: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        283: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        284: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        285: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        286: begin
          delete_size_460 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_461 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_463 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_466 <= stuckData_stuckData_3_result_0;
          delete_Key_1_467 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_470 <= stuckData_stuckData_3_result_1;
          delete_Key_2_471 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_474 <= stuckData_stuckData_3_result_2;
          delete_Key_3_475 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_478 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        287: begin
          if (delete_isLeaf_434 == 0) begin
            delete_pc <= 315;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        288: begin
          if (delete_isLeaf_461 == 0) begin
            delete_pc <= 314;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        289: begin
          delete_MergeSuccess_458 <= 0;
          case (delete_size_433)
            0: begin
              case (delete_size_460)
                0: begin
                  delete_size_433 <= delete_size_433 + 0;
                  delete_MergeSuccess_458 <= 1;
                end
                1: begin
                  delete_Key_0_436 <= delete_Key_0_463;
                  delete_Data_0_439 <= delete_Data_0_466;
                  delete_size_433 <= delete_size_433 + 1;
                  delete_MergeSuccess_458 <= 1;
                end
                2: begin
                  delete_Key_0_436 <= delete_Key_0_463;
                  delete_Data_0_439 <= delete_Data_0_466;
                  delete_Key_1_440 <= delete_Key_1_467;
                  delete_Data_1_443 <= delete_Data_1_470;
                  delete_size_433 <= delete_size_433 + 2;
                  delete_MergeSuccess_458 <= 1;
                end
                3: begin
                  delete_Key_0_436 <= delete_Key_0_463;
                  delete_Data_0_439 <= delete_Data_0_466;
                  delete_Key_1_440 <= delete_Key_1_467;
                  delete_Data_1_443 <= delete_Data_1_470;
                  delete_Key_2_444 <= delete_Key_2_471;
                  delete_Data_2_447 <= delete_Data_2_474;
                  delete_size_433 <= delete_size_433 + 3;
                  delete_MergeSuccess_458 <= 1;
                end
                4: begin
                  delete_Key_0_436 <= delete_Key_0_463;
                  delete_Data_0_439 <= delete_Data_0_466;
                  delete_Key_1_440 <= delete_Key_1_467;
                  delete_Data_1_443 <= delete_Data_1_470;
                  delete_Key_2_444 <= delete_Key_2_471;
                  delete_Data_2_447 <= delete_Data_2_474;
                  delete_Key_3_448 <= delete_Key_3_475;
                  delete_Data_3_451 <= delete_Data_3_478;
                  delete_size_433 <= delete_size_433 + 4;
                  delete_MergeSuccess_458 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_460)
                0: begin
                  delete_size_433 <= delete_size_433 + 0;
                  delete_MergeSuccess_458 <= 1;
                end
                1: begin
                  delete_Key_1_440 <= delete_Key_0_463;
                  delete_Data_1_443 <= delete_Data_0_466;
                  delete_size_433 <= delete_size_433 + 1;
                  delete_MergeSuccess_458 <= 1;
                end
                2: begin
                  delete_Key_1_440 <= delete_Key_0_463;
                  delete_Data_1_443 <= delete_Data_0_466;
                  delete_Key_2_444 <= delete_Key_1_467;
                  delete_Data_2_447 <= delete_Data_1_470;
                  delete_size_433 <= delete_size_433 + 2;
                  delete_MergeSuccess_458 <= 1;
                end
                3: begin
                  delete_Key_1_440 <= delete_Key_0_463;
                  delete_Data_1_443 <= delete_Data_0_466;
                  delete_Key_2_444 <= delete_Key_1_467;
                  delete_Data_2_447 <= delete_Data_1_470;
                  delete_Key_3_448 <= delete_Key_2_471;
                  delete_Data_3_451 <= delete_Data_2_474;
                  delete_size_433 <= delete_size_433 + 3;
                  delete_MergeSuccess_458 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_460)
                0: begin
                  delete_size_433 <= delete_size_433 + 0;
                  delete_MergeSuccess_458 <= 1;
                end
                1: begin
                  delete_Key_2_444 <= delete_Key_0_463;
                  delete_Data_2_447 <= delete_Data_0_466;
                  delete_size_433 <= delete_size_433 + 1;
                  delete_MergeSuccess_458 <= 1;
                end
                2: begin
                  delete_Key_2_444 <= delete_Key_0_463;
                  delete_Data_2_447 <= delete_Data_0_466;
                  delete_Key_3_448 <= delete_Key_1_467;
                  delete_Data_3_451 <= delete_Data_1_470;
                  delete_size_433 <= delete_size_433 + 2;
                  delete_MergeSuccess_458 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_460)
                0: begin
                  delete_size_433 <= delete_size_433 + 0;
                  delete_MergeSuccess_458 <= 1;
                end
                1: begin
                  delete_Key_3_448 <= delete_Key_0_463;
                  delete_Data_3_451 <= delete_Data_0_466;
                  delete_size_433 <= delete_size_433 + 1;
                  delete_MergeSuccess_458 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_460)
                0: begin
                  delete_size_433 <= delete_size_433 + 0;
                  delete_MergeSuccess_458 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        290: begin
          if (delete_MergeSuccess_458 == 0) begin
            delete_pc <= 313;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        291: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        292: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        293: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_488;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_488;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_488;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_488;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        294: begin
          delete_success_491 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        295: begin
          delete_stuckSize_6_index_33 <= delete_index_432;
          delete_stuckSize_6_value_34 <= delete_size_433;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_432;
          delete_stuckKeys_2_value_22 <= delete_Key_0_436;
          delete_stuckKeys_2_value_23 <= delete_Key_1_440;
          delete_stuckKeys_2_value_24 <= delete_Key_2_444;
          delete_stuckKeys_2_value_25 <= delete_Key_3_448;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_432;
          delete_stuckData_4_value_28 <= delete_Data_0_439;
          delete_stuckData_4_value_29 <= delete_Data_1_443;
          delete_stuckData_4_value_30 <= delete_Data_2_447;
          delete_stuckData_4_value_31 <= delete_Data_3_451;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        296: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        297: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        298: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        299: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        300: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        301: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        302: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        303: begin
          delete_root_494 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        304: begin
          delete_freeNext_9_index_196 <= delete_root_494;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        305: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        306: begin
          delete_next_493 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_494;
          delete_freeNext_10_value_198 <= delete_indexRight_489;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_495 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        307: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_489;
          delete_stuckIsFree_11_value_200 <= delete_isFree_495;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        308: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        309: begin
          delete_freeNext_10_index_197 <= delete_indexRight_489;
          delete_freeNext_10_value_198 <= delete_next_493;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        310: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        311: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        312: begin
          delete_pc <= 313;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        313: begin
          delete_pc <= 314;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        314: begin
          delete_pc <= 315;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        315: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 362;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        316: begin
          delete_success_557 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        317: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_554 <= delete_Data_0_82;
              delete_indexRight_555 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_554 <= delete_Data_1_86;
              delete_indexRight_555 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_554 <= delete_Data_2_90;
              delete_indexRight_555 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        318: begin
          delete_index_496 <= delete_indexLeft_554;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        319: begin
          delete_stuckSize_5_index_32 <= delete_index_496;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_496;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_496;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_496;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        320: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        321: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        322: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        323: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        324: begin
          delete_size_497 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_498 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_500 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_503 <= stuckData_stuckData_3_result_0;
          delete_Key_1_504 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_507 <= stuckData_stuckData_3_result_1;
          delete_Key_2_508 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_511 <= stuckData_stuckData_3_result_2;
          delete_Key_3_512 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_515 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        325: begin
          delete_index_523 <= delete_indexRight_555;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        326: begin
          delete_stuckSize_5_index_32 <= delete_index_523;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_523;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_523;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_523;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        327: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        328: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        329: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        330: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        331: begin
          delete_size_524 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_525 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_527 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_530 <= stuckData_stuckData_3_result_0;
          delete_Key_1_531 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_534 <= stuckData_stuckData_3_result_1;
          delete_Key_2_535 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_538 <= stuckData_stuckData_3_result_2;
          delete_Key_3_539 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_542 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        332: begin
          if (delete_isLeaf_498 == 0) begin
            delete_pc <= 334;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        333: begin
          delete_pc <= 362;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        334: begin
          if (delete_isLeaf_525 == 0) begin
            delete_pc <= 336;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        335: begin
          delete_pc <= 362;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        336: begin
          case (delete_index1_104)
            0: begin
              delete_midKey_556 <= delete_Key_0_79;
            end
            1: begin
              delete_midKey_556 <= delete_Key_1_83;
            end
            2: begin
              delete_midKey_556 <= delete_Key_2_87;
            end
            3: begin
              delete_midKey_556 <= delete_Key_3_91;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        337: begin
          delete_MergeSuccess_522 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        338: begin
          case (delete_size_497)
            0: begin
              case (delete_size_524)
                0: begin
                  delete_Key_0_500 <= delete_midKey_556;
                  delete_Data_1_507 <= delete_Data_0_530;
                  delete_size_497 <= delete_size_497 + 1;
                  delete_MergeSuccess_522 <= 1;
                end
                1: begin
                  delete_Key_0_500 <= delete_midKey_556;
                  delete_Key_1_504 <= delete_Key_0_527;
                  delete_Data_1_507 <= delete_Data_0_530;
                  delete_Data_2_511 <= delete_Data_1_534;
                  delete_size_497 <= delete_size_497 + 2;
                  delete_MergeSuccess_522 <= 1;
                end
                2: begin
                  delete_Key_0_500 <= delete_midKey_556;
                  delete_Key_1_504 <= delete_Key_0_527;
                  delete_Data_1_507 <= delete_Data_0_530;
                  delete_Key_2_508 <= delete_Key_1_531;
                  delete_Data_2_511 <= delete_Data_1_534;
                  delete_Data_3_515 <= delete_Data_2_538;
                  delete_size_497 <= delete_size_497 + 3;
                  delete_MergeSuccess_522 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_524)
                0: begin
                  delete_Key_1_504 <= delete_midKey_556;
                  delete_Data_2_511 <= delete_Data_0_530;
                  delete_size_497 <= delete_size_497 + 1;
                  delete_MergeSuccess_522 <= 1;
                end
                1: begin
                  delete_Key_1_504 <= delete_midKey_556;
                  delete_Key_2_508 <= delete_Key_0_527;
                  delete_Data_2_511 <= delete_Data_0_530;
                  delete_Data_3_515 <= delete_Data_1_534;
                  delete_size_497 <= delete_size_497 + 2;
                  delete_MergeSuccess_522 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_524)
                0: begin
                  delete_Key_2_508 <= delete_midKey_556;
                  delete_Data_3_515 <= delete_Data_0_530;
                  delete_size_497 <= delete_size_497 + 1;
                  delete_MergeSuccess_522 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_524)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_524)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        339: begin
          if (delete_MergeSuccess_522 == 0) begin
            delete_pc <= 362;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        340: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        341: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        342: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_554;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_554;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_554;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_554;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        343: begin
          delete_success_557 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        344: begin
          delete_stuckSize_6_index_33 <= delete_index_496;
          delete_stuckSize_6_value_34 <= delete_size_497;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_496;
          delete_stuckKeys_2_value_22 <= delete_Key_0_500;
          delete_stuckKeys_2_value_23 <= delete_Key_1_504;
          delete_stuckKeys_2_value_24 <= delete_Key_2_508;
          delete_stuckKeys_2_value_25 <= delete_Key_3_512;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_496;
          delete_stuckData_4_value_28 <= delete_Data_0_503;
          delete_stuckData_4_value_29 <= delete_Data_1_507;
          delete_stuckData_4_value_30 <= delete_Data_2_511;
          delete_stuckData_4_value_31 <= delete_Data_3_515;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        345: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        346: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        347: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        348: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        349: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        350: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        351: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        352: begin
          delete_root_560 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        353: begin
          delete_freeNext_9_index_196 <= delete_root_560;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        354: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        355: begin
          delete_next_559 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_560;
          delete_freeNext_10_value_198 <= delete_indexRight_555;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_561 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        356: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_555;
          delete_stuckIsFree_11_value_200 <= delete_isFree_561;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        357: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        358: begin
          delete_freeNext_10_index_197 <= delete_indexRight_555;
          delete_freeNext_10_value_198 <= delete_next_559;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        359: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        360: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        361: begin
          delete_pc <= 362;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        362: begin
          delete_pc <= 363;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2471:<init>|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        363: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 407;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        364: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_indexLeft_618 <= delete_Data_0_82;
              delete_indexRight_619 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_618 <= delete_Data_1_86;
              delete_indexRight_619 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_618 <= delete_Data_2_90;
              delete_indexRight_619 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        365: begin
          delete_index_562 <= delete_indexLeft_618;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        366: begin
          delete_stuckSize_5_index_32 <= delete_index_562;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_562;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_562;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_562;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        367: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        368: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        369: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        370: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        371: begin
          delete_size_563 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_564 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_566 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_569 <= stuckData_stuckData_3_result_0;
          delete_Key_1_570 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_573 <= stuckData_stuckData_3_result_1;
          delete_Key_2_574 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_577 <= stuckData_stuckData_3_result_2;
          delete_Key_3_578 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_581 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        372: begin
          delete_index_589 <= delete_indexRight_619;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        373: begin
          delete_stuckSize_5_index_32 <= delete_index_589;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_589;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_589;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_589;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        374: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        375: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        376: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        377: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        378: begin
          delete_size_590 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_591 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_593 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_596 <= stuckData_stuckData_3_result_0;
          delete_Key_1_597 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_600 <= stuckData_stuckData_3_result_1;
          delete_Key_2_601 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_604 <= stuckData_stuckData_3_result_2;
          delete_Key_3_605 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_608 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        379: begin
          if (delete_isLeaf_564 == 0) begin
            delete_pc <= 407;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        380: begin
          if (delete_isLeaf_591 == 0) begin
            delete_pc <= 406;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        381: begin
          delete_MergeSuccess_588 <= 0;
          case (delete_size_563)
            0: begin
              case (delete_size_590)
                0: begin
                  delete_size_563 <= delete_size_563 + 0;
                  delete_MergeSuccess_588 <= 1;
                end
                1: begin
                  delete_Key_0_566 <= delete_Key_0_593;
                  delete_Data_0_569 <= delete_Data_0_596;
                  delete_size_563 <= delete_size_563 + 1;
                  delete_MergeSuccess_588 <= 1;
                end
                2: begin
                  delete_Key_0_566 <= delete_Key_0_593;
                  delete_Data_0_569 <= delete_Data_0_596;
                  delete_Key_1_570 <= delete_Key_1_597;
                  delete_Data_1_573 <= delete_Data_1_600;
                  delete_size_563 <= delete_size_563 + 2;
                  delete_MergeSuccess_588 <= 1;
                end
                3: begin
                  delete_Key_0_566 <= delete_Key_0_593;
                  delete_Data_0_569 <= delete_Data_0_596;
                  delete_Key_1_570 <= delete_Key_1_597;
                  delete_Data_1_573 <= delete_Data_1_600;
                  delete_Key_2_574 <= delete_Key_2_601;
                  delete_Data_2_577 <= delete_Data_2_604;
                  delete_size_563 <= delete_size_563 + 3;
                  delete_MergeSuccess_588 <= 1;
                end
                4: begin
                  delete_Key_0_566 <= delete_Key_0_593;
                  delete_Data_0_569 <= delete_Data_0_596;
                  delete_Key_1_570 <= delete_Key_1_597;
                  delete_Data_1_573 <= delete_Data_1_600;
                  delete_Key_2_574 <= delete_Key_2_601;
                  delete_Data_2_577 <= delete_Data_2_604;
                  delete_Key_3_578 <= delete_Key_3_605;
                  delete_Data_3_581 <= delete_Data_3_608;
                  delete_size_563 <= delete_size_563 + 4;
                  delete_MergeSuccess_588 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_590)
                0: begin
                  delete_size_563 <= delete_size_563 + 0;
                  delete_MergeSuccess_588 <= 1;
                end
                1: begin
                  delete_Key_1_570 <= delete_Key_0_593;
                  delete_Data_1_573 <= delete_Data_0_596;
                  delete_size_563 <= delete_size_563 + 1;
                  delete_MergeSuccess_588 <= 1;
                end
                2: begin
                  delete_Key_1_570 <= delete_Key_0_593;
                  delete_Data_1_573 <= delete_Data_0_596;
                  delete_Key_2_574 <= delete_Key_1_597;
                  delete_Data_2_577 <= delete_Data_1_600;
                  delete_size_563 <= delete_size_563 + 2;
                  delete_MergeSuccess_588 <= 1;
                end
                3: begin
                  delete_Key_1_570 <= delete_Key_0_593;
                  delete_Data_1_573 <= delete_Data_0_596;
                  delete_Key_2_574 <= delete_Key_1_597;
                  delete_Data_2_577 <= delete_Data_1_600;
                  delete_Key_3_578 <= delete_Key_2_601;
                  delete_Data_3_581 <= delete_Data_2_604;
                  delete_size_563 <= delete_size_563 + 3;
                  delete_MergeSuccess_588 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_590)
                0: begin
                  delete_size_563 <= delete_size_563 + 0;
                  delete_MergeSuccess_588 <= 1;
                end
                1: begin
                  delete_Key_2_574 <= delete_Key_0_593;
                  delete_Data_2_577 <= delete_Data_0_596;
                  delete_size_563 <= delete_size_563 + 1;
                  delete_MergeSuccess_588 <= 1;
                end
                2: begin
                  delete_Key_2_574 <= delete_Key_0_593;
                  delete_Data_2_577 <= delete_Data_0_596;
                  delete_Key_3_578 <= delete_Key_1_597;
                  delete_Data_3_581 <= delete_Data_1_600;
                  delete_size_563 <= delete_size_563 + 2;
                  delete_MergeSuccess_588 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_590)
                0: begin
                  delete_size_563 <= delete_size_563 + 0;
                  delete_MergeSuccess_588 <= 1;
                end
                1: begin
                  delete_Key_3_578 <= delete_Key_0_593;
                  delete_Data_3_581 <= delete_Data_0_596;
                  delete_size_563 <= delete_size_563 + 1;
                  delete_MergeSuccess_588 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_590)
                0: begin
                  delete_size_563 <= delete_size_563 + 0;
                  delete_MergeSuccess_588 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        382: begin
          if (delete_MergeSuccess_588 == 0) begin
            delete_pc <= 405;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        383: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_StuckIndex_100) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_StuckIndex_100) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_StuckIndex_100) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        384: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        385: begin
          if (delete_StuckIndex_100 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_618;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_618;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_618;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_618;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        386: begin
          delete_success_621 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        387: begin
          delete_stuckSize_6_index_33 <= delete_index_562;
          delete_stuckSize_6_value_34 <= delete_size_563;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_562;
          delete_stuckKeys_2_value_22 <= delete_Key_0_566;
          delete_stuckKeys_2_value_23 <= delete_Key_1_570;
          delete_stuckKeys_2_value_24 <= delete_Key_2_574;
          delete_stuckKeys_2_value_25 <= delete_Key_3_578;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_562;
          delete_stuckData_4_value_28 <= delete_Data_0_569;
          delete_stuckData_4_value_29 <= delete_Data_1_573;
          delete_stuckData_4_value_30 <= delete_Data_2_577;
          delete_stuckData_4_value_31 <= delete_Data_3_581;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        388: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        389: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        390: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        391: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        392: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        393: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        394: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        395: begin
          delete_root_624 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        396: begin
          delete_freeNext_9_index_196 <= delete_root_624;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        397: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        398: begin
          delete_next_623 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_624;
          delete_freeNext_10_value_198 <= delete_indexRight_619;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_625 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        399: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_619;
          delete_stuckIsFree_11_value_200 <= delete_isFree_625;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        400: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        401: begin
          delete_freeNext_10_index_197 <= delete_indexRight_619;
          delete_freeNext_10_value_198 <= delete_next_623;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        402: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        403: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        404: begin
          delete_pc <= 405;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        405: begin
          delete_pc <= 406;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        406: begin
          delete_pc <= 407;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2476:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        407: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 454;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        408: begin
          delete_success_687 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        409: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_indexLeft_684 <= delete_Data_0_82;
              delete_indexRight_685 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_684 <= delete_Data_1_86;
              delete_indexRight_685 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_684 <= delete_Data_2_90;
              delete_indexRight_685 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        410: begin
          delete_index_626 <= delete_indexLeft_684;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        411: begin
          delete_stuckSize_5_index_32 <= delete_index_626;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_626;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_626;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_626;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        412: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        413: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        414: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        415: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        416: begin
          delete_size_627 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_628 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_630 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_633 <= stuckData_stuckData_3_result_0;
          delete_Key_1_634 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_637 <= stuckData_stuckData_3_result_1;
          delete_Key_2_638 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_641 <= stuckData_stuckData_3_result_2;
          delete_Key_3_642 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_645 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        417: begin
          delete_index_653 <= delete_indexRight_685;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        418: begin
          delete_stuckSize_5_index_32 <= delete_index_653;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_653;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_653;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_653;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        419: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        420: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        421: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        422: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        423: begin
          delete_size_654 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_655 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_657 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_660 <= stuckData_stuckData_3_result_0;
          delete_Key_1_661 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_664 <= stuckData_stuckData_3_result_1;
          delete_Key_2_665 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_668 <= stuckData_stuckData_3_result_2;
          delete_Key_3_669 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_672 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        424: begin
          if (delete_isLeaf_628 == 0) begin
            delete_pc <= 426;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        425: begin
          delete_pc <= 454;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        426: begin
          if (delete_isLeaf_655 == 0) begin
            delete_pc <= 428;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        427: begin
          delete_pc <= 454;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        428: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_midKey_686 <= delete_Key_0_79;
            end
            1: begin
              delete_midKey_686 <= delete_Key_1_83;
            end
            2: begin
              delete_midKey_686 <= delete_Key_2_87;
            end
            3: begin
              delete_midKey_686 <= delete_Key_3_91;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        429: begin
          delete_MergeSuccess_652 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        430: begin
          case (delete_size_627)
            0: begin
              case (delete_size_654)
                0: begin
                  delete_Key_0_630 <= delete_midKey_686;
                  delete_Data_1_637 <= delete_Data_0_660;
                  delete_size_627 <= delete_size_627 + 1;
                  delete_MergeSuccess_652 <= 1;
                end
                1: begin
                  delete_Key_0_630 <= delete_midKey_686;
                  delete_Key_1_634 <= delete_Key_0_657;
                  delete_Data_1_637 <= delete_Data_0_660;
                  delete_Data_2_641 <= delete_Data_1_664;
                  delete_size_627 <= delete_size_627 + 2;
                  delete_MergeSuccess_652 <= 1;
                end
                2: begin
                  delete_Key_0_630 <= delete_midKey_686;
                  delete_Key_1_634 <= delete_Key_0_657;
                  delete_Data_1_637 <= delete_Data_0_660;
                  delete_Key_2_638 <= delete_Key_1_661;
                  delete_Data_2_641 <= delete_Data_1_664;
                  delete_Data_3_645 <= delete_Data_2_668;
                  delete_size_627 <= delete_size_627 + 3;
                  delete_MergeSuccess_652 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_654)
                0: begin
                  delete_Key_1_634 <= delete_midKey_686;
                  delete_Data_2_641 <= delete_Data_0_660;
                  delete_size_627 <= delete_size_627 + 1;
                  delete_MergeSuccess_652 <= 1;
                end
                1: begin
                  delete_Key_1_634 <= delete_midKey_686;
                  delete_Key_2_638 <= delete_Key_0_657;
                  delete_Data_2_641 <= delete_Data_0_660;
                  delete_Data_3_645 <= delete_Data_1_664;
                  delete_size_627 <= delete_size_627 + 2;
                  delete_MergeSuccess_652 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_654)
                0: begin
                  delete_Key_2_638 <= delete_midKey_686;
                  delete_Data_3_645 <= delete_Data_0_660;
                  delete_size_627 <= delete_size_627 + 1;
                  delete_MergeSuccess_652 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_654)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_654)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        431: begin
          if (delete_MergeSuccess_652 == 0) begin
            delete_pc <= 454;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        432: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_StuckIndex_100) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_StuckIndex_100) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_StuckIndex_100) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        433: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        434: begin
          if (delete_StuckIndex_100 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_684;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_684;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_684;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_684;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        435: begin
          delete_success_687 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        436: begin
          delete_stuckSize_6_index_33 <= delete_index_626;
          delete_stuckSize_6_value_34 <= delete_size_627;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_626;
          delete_stuckKeys_2_value_22 <= delete_Key_0_630;
          delete_stuckKeys_2_value_23 <= delete_Key_1_634;
          delete_stuckKeys_2_value_24 <= delete_Key_2_638;
          delete_stuckKeys_2_value_25 <= delete_Key_3_642;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_626;
          delete_stuckData_4_value_28 <= delete_Data_0_633;
          delete_stuckData_4_value_29 <= delete_Data_1_637;
          delete_stuckData_4_value_30 <= delete_Data_2_641;
          delete_stuckData_4_value_31 <= delete_Data_3_645;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        437: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        438: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        439: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        440: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        441: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        442: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        443: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        444: begin
          delete_root_690 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        445: begin
          delete_freeNext_9_index_196 <= delete_root_690;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        446: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        447: begin
          delete_next_689 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_690;
          delete_freeNext_10_value_198 <= delete_indexRight_685;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_691 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        448: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_685;
          delete_stuckIsFree_11_value_200 <= delete_isFree_691;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        449: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        450: begin
          delete_freeNext_10_index_197 <= delete_indexRight_685;
          delete_freeNext_10_value_198 <= delete_next_689;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        451: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        452: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        453: begin
          delete_pc <= 454;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2477:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        454: begin
          delete_index1_104 <= delete_StuckIndex_100;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2479:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        455: begin
          delete_index1_104 <= delete_index1_104-1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0813:<init>|  Chip.java:0812:Dec|  Btree.java:2480:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        456: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 500;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        457: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_748 <= delete_Data_0_82;
              delete_indexRight_749 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_748 <= delete_Data_1_86;
              delete_indexRight_749 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_748 <= delete_Data_2_90;
              delete_indexRight_749 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        458: begin
          delete_index_692 <= delete_indexLeft_748;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        459: begin
          delete_stuckSize_5_index_32 <= delete_index_692;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_692;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_692;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_692;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        460: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        461: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        462: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        463: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        464: begin
          delete_size_693 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_694 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_696 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_699 <= stuckData_stuckData_3_result_0;
          delete_Key_1_700 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_703 <= stuckData_stuckData_3_result_1;
          delete_Key_2_704 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_707 <= stuckData_stuckData_3_result_2;
          delete_Key_3_708 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_711 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        465: begin
          delete_index_719 <= delete_indexRight_749;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        466: begin
          delete_stuckSize_5_index_32 <= delete_index_719;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_719;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_719;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_719;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        467: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        468: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        469: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        470: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        471: begin
          delete_size_720 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_721 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_723 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_726 <= stuckData_stuckData_3_result_0;
          delete_Key_1_727 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_730 <= stuckData_stuckData_3_result_1;
          delete_Key_2_731 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_734 <= stuckData_stuckData_3_result_2;
          delete_Key_3_735 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_738 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        472: begin
          if (delete_isLeaf_694 == 0) begin
            delete_pc <= 500;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        473: begin
          if (delete_isLeaf_721 == 0) begin
            delete_pc <= 499;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        474: begin
          delete_MergeSuccess_718 <= 0;
          case (delete_size_693)
            0: begin
              case (delete_size_720)
                0: begin
                  delete_size_693 <= delete_size_693 + 0;
                  delete_MergeSuccess_718 <= 1;
                end
                1: begin
                  delete_Key_0_696 <= delete_Key_0_723;
                  delete_Data_0_699 <= delete_Data_0_726;
                  delete_size_693 <= delete_size_693 + 1;
                  delete_MergeSuccess_718 <= 1;
                end
                2: begin
                  delete_Key_0_696 <= delete_Key_0_723;
                  delete_Data_0_699 <= delete_Data_0_726;
                  delete_Key_1_700 <= delete_Key_1_727;
                  delete_Data_1_703 <= delete_Data_1_730;
                  delete_size_693 <= delete_size_693 + 2;
                  delete_MergeSuccess_718 <= 1;
                end
                3: begin
                  delete_Key_0_696 <= delete_Key_0_723;
                  delete_Data_0_699 <= delete_Data_0_726;
                  delete_Key_1_700 <= delete_Key_1_727;
                  delete_Data_1_703 <= delete_Data_1_730;
                  delete_Key_2_704 <= delete_Key_2_731;
                  delete_Data_2_707 <= delete_Data_2_734;
                  delete_size_693 <= delete_size_693 + 3;
                  delete_MergeSuccess_718 <= 1;
                end
                4: begin
                  delete_Key_0_696 <= delete_Key_0_723;
                  delete_Data_0_699 <= delete_Data_0_726;
                  delete_Key_1_700 <= delete_Key_1_727;
                  delete_Data_1_703 <= delete_Data_1_730;
                  delete_Key_2_704 <= delete_Key_2_731;
                  delete_Data_2_707 <= delete_Data_2_734;
                  delete_Key_3_708 <= delete_Key_3_735;
                  delete_Data_3_711 <= delete_Data_3_738;
                  delete_size_693 <= delete_size_693 + 4;
                  delete_MergeSuccess_718 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_720)
                0: begin
                  delete_size_693 <= delete_size_693 + 0;
                  delete_MergeSuccess_718 <= 1;
                end
                1: begin
                  delete_Key_1_700 <= delete_Key_0_723;
                  delete_Data_1_703 <= delete_Data_0_726;
                  delete_size_693 <= delete_size_693 + 1;
                  delete_MergeSuccess_718 <= 1;
                end
                2: begin
                  delete_Key_1_700 <= delete_Key_0_723;
                  delete_Data_1_703 <= delete_Data_0_726;
                  delete_Key_2_704 <= delete_Key_1_727;
                  delete_Data_2_707 <= delete_Data_1_730;
                  delete_size_693 <= delete_size_693 + 2;
                  delete_MergeSuccess_718 <= 1;
                end
                3: begin
                  delete_Key_1_700 <= delete_Key_0_723;
                  delete_Data_1_703 <= delete_Data_0_726;
                  delete_Key_2_704 <= delete_Key_1_727;
                  delete_Data_2_707 <= delete_Data_1_730;
                  delete_Key_3_708 <= delete_Key_2_731;
                  delete_Data_3_711 <= delete_Data_2_734;
                  delete_size_693 <= delete_size_693 + 3;
                  delete_MergeSuccess_718 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_720)
                0: begin
                  delete_size_693 <= delete_size_693 + 0;
                  delete_MergeSuccess_718 <= 1;
                end
                1: begin
                  delete_Key_2_704 <= delete_Key_0_723;
                  delete_Data_2_707 <= delete_Data_0_726;
                  delete_size_693 <= delete_size_693 + 1;
                  delete_MergeSuccess_718 <= 1;
                end
                2: begin
                  delete_Key_2_704 <= delete_Key_0_723;
                  delete_Data_2_707 <= delete_Data_0_726;
                  delete_Key_3_708 <= delete_Key_1_727;
                  delete_Data_3_711 <= delete_Data_1_730;
                  delete_size_693 <= delete_size_693 + 2;
                  delete_MergeSuccess_718 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_720)
                0: begin
                  delete_size_693 <= delete_size_693 + 0;
                  delete_MergeSuccess_718 <= 1;
                end
                1: begin
                  delete_Key_3_708 <= delete_Key_0_723;
                  delete_Data_3_711 <= delete_Data_0_726;
                  delete_size_693 <= delete_size_693 + 1;
                  delete_MergeSuccess_718 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_720)
                0: begin
                  delete_size_693 <= delete_size_693 + 0;
                  delete_MergeSuccess_718 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        475: begin
          if (delete_MergeSuccess_718 == 0) begin
            delete_pc <= 498;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        476: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        477: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        478: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_748;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_748;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_748;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_748;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        479: begin
          delete_success_751 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        480: begin
          delete_stuckSize_6_index_33 <= delete_index_692;
          delete_stuckSize_6_value_34 <= delete_size_693;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_692;
          delete_stuckKeys_2_value_22 <= delete_Key_0_696;
          delete_stuckKeys_2_value_23 <= delete_Key_1_700;
          delete_stuckKeys_2_value_24 <= delete_Key_2_704;
          delete_stuckKeys_2_value_25 <= delete_Key_3_708;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_692;
          delete_stuckData_4_value_28 <= delete_Data_0_699;
          delete_stuckData_4_value_29 <= delete_Data_1_703;
          delete_stuckData_4_value_30 <= delete_Data_2_707;
          delete_stuckData_4_value_31 <= delete_Data_3_711;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        481: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        482: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        483: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        484: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        485: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        486: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        487: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        488: begin
          delete_root_754 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        489: begin
          delete_freeNext_9_index_196 <= delete_root_754;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        490: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        491: begin
          delete_next_753 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_754;
          delete_freeNext_10_value_198 <= delete_indexRight_749;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_755 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        492: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_749;
          delete_stuckIsFree_11_value_200 <= delete_isFree_755;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        493: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        494: begin
          delete_freeNext_10_index_197 <= delete_indexRight_749;
          delete_freeNext_10_value_198 <= delete_next_753;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        495: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        496: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        497: begin
          delete_pc <= 498;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        498: begin
          delete_pc <= 499;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        499: begin
          delete_pc <= 500;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2481:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        500: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 547;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        501: begin
          delete_success_817 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        502: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_814 <= delete_Data_0_82;
              delete_indexRight_815 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_814 <= delete_Data_1_86;
              delete_indexRight_815 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_814 <= delete_Data_2_90;
              delete_indexRight_815 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        503: begin
          delete_index_756 <= delete_indexLeft_814;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        504: begin
          delete_stuckSize_5_index_32 <= delete_index_756;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_756;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_756;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_756;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        505: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        506: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        507: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        508: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        509: begin
          delete_size_757 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_758 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_760 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_763 <= stuckData_stuckData_3_result_0;
          delete_Key_1_764 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_767 <= stuckData_stuckData_3_result_1;
          delete_Key_2_768 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_771 <= stuckData_stuckData_3_result_2;
          delete_Key_3_772 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_775 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        510: begin
          delete_index_783 <= delete_indexRight_815;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        511: begin
          delete_stuckSize_5_index_32 <= delete_index_783;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_783;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_783;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_783;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        512: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        513: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        514: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        515: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        516: begin
          delete_size_784 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_785 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_787 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_790 <= stuckData_stuckData_3_result_0;
          delete_Key_1_791 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_794 <= stuckData_stuckData_3_result_1;
          delete_Key_2_795 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_798 <= stuckData_stuckData_3_result_2;
          delete_Key_3_799 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_802 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        517: begin
          if (delete_isLeaf_758 == 0) begin
            delete_pc <= 519;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        518: begin
          delete_pc <= 547;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        519: begin
          if (delete_isLeaf_785 == 0) begin
            delete_pc <= 521;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        520: begin
          delete_pc <= 547;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        521: begin
          case (delete_index1_104)
            0: begin
              delete_midKey_816 <= delete_Key_0_79;
            end
            1: begin
              delete_midKey_816 <= delete_Key_1_83;
            end
            2: begin
              delete_midKey_816 <= delete_Key_2_87;
            end
            3: begin
              delete_midKey_816 <= delete_Key_3_91;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        522: begin
          delete_MergeSuccess_782 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        523: begin
          case (delete_size_757)
            0: begin
              case (delete_size_784)
                0: begin
                  delete_Key_0_760 <= delete_midKey_816;
                  delete_Data_1_767 <= delete_Data_0_790;
                  delete_size_757 <= delete_size_757 + 1;
                  delete_MergeSuccess_782 <= 1;
                end
                1: begin
                  delete_Key_0_760 <= delete_midKey_816;
                  delete_Key_1_764 <= delete_Key_0_787;
                  delete_Data_1_767 <= delete_Data_0_790;
                  delete_Data_2_771 <= delete_Data_1_794;
                  delete_size_757 <= delete_size_757 + 2;
                  delete_MergeSuccess_782 <= 1;
                end
                2: begin
                  delete_Key_0_760 <= delete_midKey_816;
                  delete_Key_1_764 <= delete_Key_0_787;
                  delete_Data_1_767 <= delete_Data_0_790;
                  delete_Key_2_768 <= delete_Key_1_791;
                  delete_Data_2_771 <= delete_Data_1_794;
                  delete_Data_3_775 <= delete_Data_2_798;
                  delete_size_757 <= delete_size_757 + 3;
                  delete_MergeSuccess_782 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_784)
                0: begin
                  delete_Key_1_764 <= delete_midKey_816;
                  delete_Data_2_771 <= delete_Data_0_790;
                  delete_size_757 <= delete_size_757 + 1;
                  delete_MergeSuccess_782 <= 1;
                end
                1: begin
                  delete_Key_1_764 <= delete_midKey_816;
                  delete_Key_2_768 <= delete_Key_0_787;
                  delete_Data_2_771 <= delete_Data_0_790;
                  delete_Data_3_775 <= delete_Data_1_794;
                  delete_size_757 <= delete_size_757 + 2;
                  delete_MergeSuccess_782 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_784)
                0: begin
                  delete_Key_2_768 <= delete_midKey_816;
                  delete_Data_3_775 <= delete_Data_0_790;
                  delete_size_757 <= delete_size_757 + 1;
                  delete_MergeSuccess_782 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_784)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_784)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        524: begin
          if (delete_MergeSuccess_782 == 0) begin
            delete_pc <= 547;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        525: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        526: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        527: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_814;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_814;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_814;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_814;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        528: begin
          delete_success_817 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        529: begin
          delete_stuckSize_6_index_33 <= delete_index_756;
          delete_stuckSize_6_value_34 <= delete_size_757;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_756;
          delete_stuckKeys_2_value_22 <= delete_Key_0_760;
          delete_stuckKeys_2_value_23 <= delete_Key_1_764;
          delete_stuckKeys_2_value_24 <= delete_Key_2_768;
          delete_stuckKeys_2_value_25 <= delete_Key_3_772;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_756;
          delete_stuckData_4_value_28 <= delete_Data_0_763;
          delete_stuckData_4_value_29 <= delete_Data_1_767;
          delete_stuckData_4_value_30 <= delete_Data_2_771;
          delete_stuckData_4_value_31 <= delete_Data_3_775;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        530: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        531: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        532: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        533: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        534: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        535: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        536: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        537: begin
          delete_root_820 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        538: begin
          delete_freeNext_9_index_196 <= delete_root_820;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        539: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        540: begin
          delete_next_819 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_820;
          delete_freeNext_10_value_198 <= delete_indexRight_815;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_821 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        541: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_815;
          delete_stuckIsFree_11_value_200 <= delete_isFree_821;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        542: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        543: begin
          delete_freeNext_10_index_197 <= delete_indexRight_815;
          delete_freeNext_10_value_198 <= delete_next_819;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        544: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        545: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        546: begin
          delete_pc <= 547;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2482:Then|  Chip.java:0610:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        547: begin
          delete_pc <= 730;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        548: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 592;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        549: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_878 <= delete_Data_0_82;
              delete_indexRight_879 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_878 <= delete_Data_1_86;
              delete_indexRight_879 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_878 <= delete_Data_2_90;
              delete_indexRight_879 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        550: begin
          delete_index_822 <= delete_indexLeft_878;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        551: begin
          delete_stuckSize_5_index_32 <= delete_index_822;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_822;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_822;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_822;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        552: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        553: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        554: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        555: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        556: begin
          delete_size_823 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_824 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_826 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_829 <= stuckData_stuckData_3_result_0;
          delete_Key_1_830 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_833 <= stuckData_stuckData_3_result_1;
          delete_Key_2_834 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_837 <= stuckData_stuckData_3_result_2;
          delete_Key_3_838 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_841 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        557: begin
          delete_index_849 <= delete_indexRight_879;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        558: begin
          delete_stuckSize_5_index_32 <= delete_index_849;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_849;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_849;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_849;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        559: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        560: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        561: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        562: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        563: begin
          delete_size_850 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_851 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_853 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_856 <= stuckData_stuckData_3_result_0;
          delete_Key_1_857 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_860 <= stuckData_stuckData_3_result_1;
          delete_Key_2_861 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_864 <= stuckData_stuckData_3_result_2;
          delete_Key_3_865 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_868 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        564: begin
          if (delete_isLeaf_824 == 0) begin
            delete_pc <= 592;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        565: begin
          if (delete_isLeaf_851 == 0) begin
            delete_pc <= 591;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        566: begin
          delete_MergeSuccess_848 <= 0;
          case (delete_size_823)
            0: begin
              case (delete_size_850)
                0: begin
                  delete_size_823 <= delete_size_823 + 0;
                  delete_MergeSuccess_848 <= 1;
                end
                1: begin
                  delete_Key_0_826 <= delete_Key_0_853;
                  delete_Data_0_829 <= delete_Data_0_856;
                  delete_size_823 <= delete_size_823 + 1;
                  delete_MergeSuccess_848 <= 1;
                end
                2: begin
                  delete_Key_0_826 <= delete_Key_0_853;
                  delete_Data_0_829 <= delete_Data_0_856;
                  delete_Key_1_830 <= delete_Key_1_857;
                  delete_Data_1_833 <= delete_Data_1_860;
                  delete_size_823 <= delete_size_823 + 2;
                  delete_MergeSuccess_848 <= 1;
                end
                3: begin
                  delete_Key_0_826 <= delete_Key_0_853;
                  delete_Data_0_829 <= delete_Data_0_856;
                  delete_Key_1_830 <= delete_Key_1_857;
                  delete_Data_1_833 <= delete_Data_1_860;
                  delete_Key_2_834 <= delete_Key_2_861;
                  delete_Data_2_837 <= delete_Data_2_864;
                  delete_size_823 <= delete_size_823 + 3;
                  delete_MergeSuccess_848 <= 1;
                end
                4: begin
                  delete_Key_0_826 <= delete_Key_0_853;
                  delete_Data_0_829 <= delete_Data_0_856;
                  delete_Key_1_830 <= delete_Key_1_857;
                  delete_Data_1_833 <= delete_Data_1_860;
                  delete_Key_2_834 <= delete_Key_2_861;
                  delete_Data_2_837 <= delete_Data_2_864;
                  delete_Key_3_838 <= delete_Key_3_865;
                  delete_Data_3_841 <= delete_Data_3_868;
                  delete_size_823 <= delete_size_823 + 4;
                  delete_MergeSuccess_848 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_850)
                0: begin
                  delete_size_823 <= delete_size_823 + 0;
                  delete_MergeSuccess_848 <= 1;
                end
                1: begin
                  delete_Key_1_830 <= delete_Key_0_853;
                  delete_Data_1_833 <= delete_Data_0_856;
                  delete_size_823 <= delete_size_823 + 1;
                  delete_MergeSuccess_848 <= 1;
                end
                2: begin
                  delete_Key_1_830 <= delete_Key_0_853;
                  delete_Data_1_833 <= delete_Data_0_856;
                  delete_Key_2_834 <= delete_Key_1_857;
                  delete_Data_2_837 <= delete_Data_1_860;
                  delete_size_823 <= delete_size_823 + 2;
                  delete_MergeSuccess_848 <= 1;
                end
                3: begin
                  delete_Key_1_830 <= delete_Key_0_853;
                  delete_Data_1_833 <= delete_Data_0_856;
                  delete_Key_2_834 <= delete_Key_1_857;
                  delete_Data_2_837 <= delete_Data_1_860;
                  delete_Key_3_838 <= delete_Key_2_861;
                  delete_Data_3_841 <= delete_Data_2_864;
                  delete_size_823 <= delete_size_823 + 3;
                  delete_MergeSuccess_848 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_850)
                0: begin
                  delete_size_823 <= delete_size_823 + 0;
                  delete_MergeSuccess_848 <= 1;
                end
                1: begin
                  delete_Key_2_834 <= delete_Key_0_853;
                  delete_Data_2_837 <= delete_Data_0_856;
                  delete_size_823 <= delete_size_823 + 1;
                  delete_MergeSuccess_848 <= 1;
                end
                2: begin
                  delete_Key_2_834 <= delete_Key_0_853;
                  delete_Data_2_837 <= delete_Data_0_856;
                  delete_Key_3_838 <= delete_Key_1_857;
                  delete_Data_3_841 <= delete_Data_1_860;
                  delete_size_823 <= delete_size_823 + 2;
                  delete_MergeSuccess_848 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_850)
                0: begin
                  delete_size_823 <= delete_size_823 + 0;
                  delete_MergeSuccess_848 <= 1;
                end
                1: begin
                  delete_Key_3_838 <= delete_Key_0_853;
                  delete_Data_3_841 <= delete_Data_0_856;
                  delete_size_823 <= delete_size_823 + 1;
                  delete_MergeSuccess_848 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_850)
                0: begin
                  delete_size_823 <= delete_size_823 + 0;
                  delete_MergeSuccess_848 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        567: begin
          if (delete_MergeSuccess_848 == 0) begin
            delete_pc <= 590;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        568: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        569: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        570: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_878;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_878;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_878;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_878;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        571: begin
          delete_success_881 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        572: begin
          delete_stuckSize_6_index_33 <= delete_index_822;
          delete_stuckSize_6_value_34 <= delete_size_823;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_822;
          delete_stuckKeys_2_value_22 <= delete_Key_0_826;
          delete_stuckKeys_2_value_23 <= delete_Key_1_830;
          delete_stuckKeys_2_value_24 <= delete_Key_2_834;
          delete_stuckKeys_2_value_25 <= delete_Key_3_838;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_822;
          delete_stuckData_4_value_28 <= delete_Data_0_829;
          delete_stuckData_4_value_29 <= delete_Data_1_833;
          delete_stuckData_4_value_30 <= delete_Data_2_837;
          delete_stuckData_4_value_31 <= delete_Data_3_841;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        573: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        574: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        575: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        576: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        577: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        578: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        579: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        580: begin
          delete_root_884 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        581: begin
          delete_freeNext_9_index_196 <= delete_root_884;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        582: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        583: begin
          delete_next_883 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_884;
          delete_freeNext_10_value_198 <= delete_indexRight_879;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_885 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        584: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_879;
          delete_stuckIsFree_11_value_200 <= delete_isFree_885;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        585: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        586: begin
          delete_freeNext_10_index_197 <= delete_indexRight_879;
          delete_freeNext_10_value_198 <= delete_next_883;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        587: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        588: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        589: begin
          delete_pc <= 590;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        590: begin
          delete_pc <= 591;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        591: begin
          delete_pc <= 592;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2486:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        592: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 639;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        593: begin
          delete_success_947 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        594: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_944 <= delete_Data_0_82;
              delete_indexRight_945 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_944 <= delete_Data_1_86;
              delete_indexRight_945 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_944 <= delete_Data_2_90;
              delete_indexRight_945 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        595: begin
          delete_index_886 <= delete_indexLeft_944;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        596: begin
          delete_stuckSize_5_index_32 <= delete_index_886;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_886;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_886;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_886;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        597: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        598: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        599: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        600: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        601: begin
          delete_size_887 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_888 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_890 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_893 <= stuckData_stuckData_3_result_0;
          delete_Key_1_894 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_897 <= stuckData_stuckData_3_result_1;
          delete_Key_2_898 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_901 <= stuckData_stuckData_3_result_2;
          delete_Key_3_902 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_905 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        602: begin
          delete_index_913 <= delete_indexRight_945;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        603: begin
          delete_stuckSize_5_index_32 <= delete_index_913;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_913;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_913;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_913;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        604: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        605: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        606: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        607: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        608: begin
          delete_size_914 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_915 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_917 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_920 <= stuckData_stuckData_3_result_0;
          delete_Key_1_921 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_924 <= stuckData_stuckData_3_result_1;
          delete_Key_2_925 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_928 <= stuckData_stuckData_3_result_2;
          delete_Key_3_929 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_932 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        609: begin
          if (delete_isLeaf_888 == 0) begin
            delete_pc <= 611;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        610: begin
          delete_pc <= 639;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        611: begin
          if (delete_isLeaf_915 == 0) begin
            delete_pc <= 613;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        612: begin
          delete_pc <= 639;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        613: begin
          case (delete_index1_104)
            0: begin
              delete_midKey_946 <= delete_Key_0_79;
            end
            1: begin
              delete_midKey_946 <= delete_Key_1_83;
            end
            2: begin
              delete_midKey_946 <= delete_Key_2_87;
            end
            3: begin
              delete_midKey_946 <= delete_Key_3_91;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        614: begin
          delete_MergeSuccess_912 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        615: begin
          case (delete_size_887)
            0: begin
              case (delete_size_914)
                0: begin
                  delete_Key_0_890 <= delete_midKey_946;
                  delete_Data_1_897 <= delete_Data_0_920;
                  delete_size_887 <= delete_size_887 + 1;
                  delete_MergeSuccess_912 <= 1;
                end
                1: begin
                  delete_Key_0_890 <= delete_midKey_946;
                  delete_Key_1_894 <= delete_Key_0_917;
                  delete_Data_1_897 <= delete_Data_0_920;
                  delete_Data_2_901 <= delete_Data_1_924;
                  delete_size_887 <= delete_size_887 + 2;
                  delete_MergeSuccess_912 <= 1;
                end
                2: begin
                  delete_Key_0_890 <= delete_midKey_946;
                  delete_Key_1_894 <= delete_Key_0_917;
                  delete_Data_1_897 <= delete_Data_0_920;
                  delete_Key_2_898 <= delete_Key_1_921;
                  delete_Data_2_901 <= delete_Data_1_924;
                  delete_Data_3_905 <= delete_Data_2_928;
                  delete_size_887 <= delete_size_887 + 3;
                  delete_MergeSuccess_912 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_914)
                0: begin
                  delete_Key_1_894 <= delete_midKey_946;
                  delete_Data_2_901 <= delete_Data_0_920;
                  delete_size_887 <= delete_size_887 + 1;
                  delete_MergeSuccess_912 <= 1;
                end
                1: begin
                  delete_Key_1_894 <= delete_midKey_946;
                  delete_Key_2_898 <= delete_Key_0_917;
                  delete_Data_2_901 <= delete_Data_0_920;
                  delete_Data_3_905 <= delete_Data_1_924;
                  delete_size_887 <= delete_size_887 + 2;
                  delete_MergeSuccess_912 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_914)
                0: begin
                  delete_Key_2_898 <= delete_midKey_946;
                  delete_Data_3_905 <= delete_Data_0_920;
                  delete_size_887 <= delete_size_887 + 1;
                  delete_MergeSuccess_912 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_914)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_914)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        616: begin
          if (delete_MergeSuccess_912 == 0) begin
            delete_pc <= 639;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        617: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        618: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        619: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_944;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_944;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_944;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_944;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        620: begin
          delete_success_947 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        621: begin
          delete_stuckSize_6_index_33 <= delete_index_886;
          delete_stuckSize_6_value_34 <= delete_size_887;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_886;
          delete_stuckKeys_2_value_22 <= delete_Key_0_890;
          delete_stuckKeys_2_value_23 <= delete_Key_1_894;
          delete_stuckKeys_2_value_24 <= delete_Key_2_898;
          delete_stuckKeys_2_value_25 <= delete_Key_3_902;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_886;
          delete_stuckData_4_value_28 <= delete_Data_0_893;
          delete_stuckData_4_value_29 <= delete_Data_1_897;
          delete_stuckData_4_value_30 <= delete_Data_2_901;
          delete_stuckData_4_value_31 <= delete_Data_3_905;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        622: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        623: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        624: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        625: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        626: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        627: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        628: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        629: begin
          delete_root_950 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        630: begin
          delete_freeNext_9_index_196 <= delete_root_950;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        631: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        632: begin
          delete_next_949 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_950;
          delete_freeNext_10_value_198 <= delete_indexRight_945;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_951 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        633: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_945;
          delete_stuckIsFree_11_value_200 <= delete_isFree_951;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        634: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        635: begin
          delete_freeNext_10_index_197 <= delete_indexRight_945;
          delete_freeNext_10_value_198 <= delete_next_949;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        636: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        637: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        638: begin
          delete_pc <= 639;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2487:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        639: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 683;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        640: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_indexLeft_1008 <= delete_Data_0_82;
              delete_indexRight_1009 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_1008 <= delete_Data_1_86;
              delete_indexRight_1009 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_1008 <= delete_Data_2_90;
              delete_indexRight_1009 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        641: begin
          delete_index_952 <= delete_indexLeft_1008;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        642: begin
          delete_stuckSize_5_index_32 <= delete_index_952;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_952;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_952;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_952;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        643: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        644: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        645: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        646: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        647: begin
          delete_size_953 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_954 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_956 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_959 <= stuckData_stuckData_3_result_0;
          delete_Key_1_960 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_963 <= stuckData_stuckData_3_result_1;
          delete_Key_2_964 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_967 <= stuckData_stuckData_3_result_2;
          delete_Key_3_968 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_971 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        648: begin
          delete_index_979 <= delete_indexRight_1009;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        649: begin
          delete_stuckSize_5_index_32 <= delete_index_979;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_979;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_979;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_979;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        650: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        651: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        652: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        653: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        654: begin
          delete_size_980 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_981 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_983 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_986 <= stuckData_stuckData_3_result_0;
          delete_Key_1_987 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_990 <= stuckData_stuckData_3_result_1;
          delete_Key_2_991 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_994 <= stuckData_stuckData_3_result_2;
          delete_Key_3_995 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_998 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        655: begin
          if (delete_isLeaf_954 == 0) begin
            delete_pc <= 683;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        656: begin
          if (delete_isLeaf_981 == 0) begin
            delete_pc <= 682;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        657: begin
          delete_MergeSuccess_978 <= 0;
          case (delete_size_953)
            0: begin
              case (delete_size_980)
                0: begin
                  delete_size_953 <= delete_size_953 + 0;
                  delete_MergeSuccess_978 <= 1;
                end
                1: begin
                  delete_Key_0_956 <= delete_Key_0_983;
                  delete_Data_0_959 <= delete_Data_0_986;
                  delete_size_953 <= delete_size_953 + 1;
                  delete_MergeSuccess_978 <= 1;
                end
                2: begin
                  delete_Key_0_956 <= delete_Key_0_983;
                  delete_Data_0_959 <= delete_Data_0_986;
                  delete_Key_1_960 <= delete_Key_1_987;
                  delete_Data_1_963 <= delete_Data_1_990;
                  delete_size_953 <= delete_size_953 + 2;
                  delete_MergeSuccess_978 <= 1;
                end
                3: begin
                  delete_Key_0_956 <= delete_Key_0_983;
                  delete_Data_0_959 <= delete_Data_0_986;
                  delete_Key_1_960 <= delete_Key_1_987;
                  delete_Data_1_963 <= delete_Data_1_990;
                  delete_Key_2_964 <= delete_Key_2_991;
                  delete_Data_2_967 <= delete_Data_2_994;
                  delete_size_953 <= delete_size_953 + 3;
                  delete_MergeSuccess_978 <= 1;
                end
                4: begin
                  delete_Key_0_956 <= delete_Key_0_983;
                  delete_Data_0_959 <= delete_Data_0_986;
                  delete_Key_1_960 <= delete_Key_1_987;
                  delete_Data_1_963 <= delete_Data_1_990;
                  delete_Key_2_964 <= delete_Key_2_991;
                  delete_Data_2_967 <= delete_Data_2_994;
                  delete_Key_3_968 <= delete_Key_3_995;
                  delete_Data_3_971 <= delete_Data_3_998;
                  delete_size_953 <= delete_size_953 + 4;
                  delete_MergeSuccess_978 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_980)
                0: begin
                  delete_size_953 <= delete_size_953 + 0;
                  delete_MergeSuccess_978 <= 1;
                end
                1: begin
                  delete_Key_1_960 <= delete_Key_0_983;
                  delete_Data_1_963 <= delete_Data_0_986;
                  delete_size_953 <= delete_size_953 + 1;
                  delete_MergeSuccess_978 <= 1;
                end
                2: begin
                  delete_Key_1_960 <= delete_Key_0_983;
                  delete_Data_1_963 <= delete_Data_0_986;
                  delete_Key_2_964 <= delete_Key_1_987;
                  delete_Data_2_967 <= delete_Data_1_990;
                  delete_size_953 <= delete_size_953 + 2;
                  delete_MergeSuccess_978 <= 1;
                end
                3: begin
                  delete_Key_1_960 <= delete_Key_0_983;
                  delete_Data_1_963 <= delete_Data_0_986;
                  delete_Key_2_964 <= delete_Key_1_987;
                  delete_Data_2_967 <= delete_Data_1_990;
                  delete_Key_3_968 <= delete_Key_2_991;
                  delete_Data_3_971 <= delete_Data_2_994;
                  delete_size_953 <= delete_size_953 + 3;
                  delete_MergeSuccess_978 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_980)
                0: begin
                  delete_size_953 <= delete_size_953 + 0;
                  delete_MergeSuccess_978 <= 1;
                end
                1: begin
                  delete_Key_2_964 <= delete_Key_0_983;
                  delete_Data_2_967 <= delete_Data_0_986;
                  delete_size_953 <= delete_size_953 + 1;
                  delete_MergeSuccess_978 <= 1;
                end
                2: begin
                  delete_Key_2_964 <= delete_Key_0_983;
                  delete_Data_2_967 <= delete_Data_0_986;
                  delete_Key_3_968 <= delete_Key_1_987;
                  delete_Data_3_971 <= delete_Data_1_990;
                  delete_size_953 <= delete_size_953 + 2;
                  delete_MergeSuccess_978 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_980)
                0: begin
                  delete_size_953 <= delete_size_953 + 0;
                  delete_MergeSuccess_978 <= 1;
                end
                1: begin
                  delete_Key_3_968 <= delete_Key_0_983;
                  delete_Data_3_971 <= delete_Data_0_986;
                  delete_size_953 <= delete_size_953 + 1;
                  delete_MergeSuccess_978 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_980)
                0: begin
                  delete_size_953 <= delete_size_953 + 0;
                  delete_MergeSuccess_978 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        658: begin
          if (delete_MergeSuccess_978 == 0) begin
            delete_pc <= 681;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        659: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_StuckIndex_100) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_StuckIndex_100) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_StuckIndex_100) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        660: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        661: begin
          if (delete_StuckIndex_100 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_1008;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_1008;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_1008;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_1008;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        662: begin
          delete_success_1011 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        663: begin
          delete_stuckSize_6_index_33 <= delete_index_952;
          delete_stuckSize_6_value_34 <= delete_size_953;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_952;
          delete_stuckKeys_2_value_22 <= delete_Key_0_956;
          delete_stuckKeys_2_value_23 <= delete_Key_1_960;
          delete_stuckKeys_2_value_24 <= delete_Key_2_964;
          delete_stuckKeys_2_value_25 <= delete_Key_3_968;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_952;
          delete_stuckData_4_value_28 <= delete_Data_0_959;
          delete_stuckData_4_value_29 <= delete_Data_1_963;
          delete_stuckData_4_value_30 <= delete_Data_2_967;
          delete_stuckData_4_value_31 <= delete_Data_3_971;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        664: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        665: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        666: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        667: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        668: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        669: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        670: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        671: begin
          delete_root_1014 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        672: begin
          delete_freeNext_9_index_196 <= delete_root_1014;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        673: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        674: begin
          delete_next_1013 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_1014;
          delete_freeNext_10_value_198 <= delete_indexRight_1009;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_1015 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        675: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_1009;
          delete_stuckIsFree_11_value_200 <= delete_isFree_1015;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        676: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        677: begin
          delete_freeNext_10_index_197 <= delete_indexRight_1009;
          delete_freeNext_10_value_198 <= delete_next_1013;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        678: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        679: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        680: begin
          delete_pc <= 681;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        681: begin
          delete_pc <= 682;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        682: begin
          delete_pc <= 683;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2489:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        683: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 730;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        684: begin
          delete_success_1077 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        685: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_indexLeft_1074 <= delete_Data_0_82;
              delete_indexRight_1075 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_1074 <= delete_Data_1_86;
              delete_indexRight_1075 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_1074 <= delete_Data_2_90;
              delete_indexRight_1075 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        686: begin
          delete_index_1016 <= delete_indexLeft_1074;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        687: begin
          delete_stuckSize_5_index_32 <= delete_index_1016;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_1016;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_1016;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_1016;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        688: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        689: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        690: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        691: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        692: begin
          delete_size_1017 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_1018 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_1020 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_1023 <= stuckData_stuckData_3_result_0;
          delete_Key_1_1024 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_1027 <= stuckData_stuckData_3_result_1;
          delete_Key_2_1028 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_1031 <= stuckData_stuckData_3_result_2;
          delete_Key_3_1032 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_1035 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        693: begin
          delete_index_1043 <= delete_indexRight_1075;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        694: begin
          delete_stuckSize_5_index_32 <= delete_index_1043;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_1043;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_1043;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_1043;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        695: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        696: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        697: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        698: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        699: begin
          delete_size_1044 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_1045 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_1047 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_1050 <= stuckData_stuckData_3_result_0;
          delete_Key_1_1051 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_1054 <= stuckData_stuckData_3_result_1;
          delete_Key_2_1055 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_1058 <= stuckData_stuckData_3_result_2;
          delete_Key_3_1059 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_1062 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        700: begin
          if (delete_isLeaf_1018 == 0) begin
            delete_pc <= 702;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        701: begin
          delete_pc <= 730;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        702: begin
          if (delete_isLeaf_1045 == 0) begin
            delete_pc <= 704;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        703: begin
          delete_pc <= 730;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        704: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_midKey_1076 <= delete_Key_0_79;
            end
            1: begin
              delete_midKey_1076 <= delete_Key_1_83;
            end
            2: begin
              delete_midKey_1076 <= delete_Key_2_87;
            end
            3: begin
              delete_midKey_1076 <= delete_Key_3_91;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        705: begin
          delete_MergeSuccess_1042 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        706: begin
          case (delete_size_1017)
            0: begin
              case (delete_size_1044)
                0: begin
                  delete_Key_0_1020 <= delete_midKey_1076;
                  delete_Data_1_1027 <= delete_Data_0_1050;
                  delete_size_1017 <= delete_size_1017 + 1;
                  delete_MergeSuccess_1042 <= 1;
                end
                1: begin
                  delete_Key_0_1020 <= delete_midKey_1076;
                  delete_Key_1_1024 <= delete_Key_0_1047;
                  delete_Data_1_1027 <= delete_Data_0_1050;
                  delete_Data_2_1031 <= delete_Data_1_1054;
                  delete_size_1017 <= delete_size_1017 + 2;
                  delete_MergeSuccess_1042 <= 1;
                end
                2: begin
                  delete_Key_0_1020 <= delete_midKey_1076;
                  delete_Key_1_1024 <= delete_Key_0_1047;
                  delete_Data_1_1027 <= delete_Data_0_1050;
                  delete_Key_2_1028 <= delete_Key_1_1051;
                  delete_Data_2_1031 <= delete_Data_1_1054;
                  delete_Data_3_1035 <= delete_Data_2_1058;
                  delete_size_1017 <= delete_size_1017 + 3;
                  delete_MergeSuccess_1042 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_1044)
                0: begin
                  delete_Key_1_1024 <= delete_midKey_1076;
                  delete_Data_2_1031 <= delete_Data_0_1050;
                  delete_size_1017 <= delete_size_1017 + 1;
                  delete_MergeSuccess_1042 <= 1;
                end
                1: begin
                  delete_Key_1_1024 <= delete_midKey_1076;
                  delete_Key_2_1028 <= delete_Key_0_1047;
                  delete_Data_2_1031 <= delete_Data_0_1050;
                  delete_Data_3_1035 <= delete_Data_1_1054;
                  delete_size_1017 <= delete_size_1017 + 2;
                  delete_MergeSuccess_1042 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_1044)
                0: begin
                  delete_Key_2_1028 <= delete_midKey_1076;
                  delete_Data_3_1035 <= delete_Data_0_1050;
                  delete_size_1017 <= delete_size_1017 + 1;
                  delete_MergeSuccess_1042 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_1044)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_1044)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        707: begin
          if (delete_MergeSuccess_1042 == 0) begin
            delete_pc <= 730;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        708: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_StuckIndex_100) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_StuckIndex_100) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_StuckIndex_100) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        709: begin
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        710: begin
          if (delete_StuckIndex_100 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_StuckIndex_100)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_1074;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_1074;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_1074;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_1074;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        711: begin
          delete_success_1077 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        712: begin
          delete_stuckSize_6_index_33 <= delete_index_1016;
          delete_stuckSize_6_value_34 <= delete_size_1017;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_1016;
          delete_stuckKeys_2_value_22 <= delete_Key_0_1020;
          delete_stuckKeys_2_value_23 <= delete_Key_1_1024;
          delete_stuckKeys_2_value_24 <= delete_Key_2_1028;
          delete_stuckKeys_2_value_25 <= delete_Key_3_1032;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_1016;
          delete_stuckData_4_value_28 <= delete_Data_0_1023;
          delete_stuckData_4_value_29 <= delete_Data_1_1027;
          delete_stuckData_4_value_30 <= delete_Data_2_1031;
          delete_stuckData_4_value_31 <= delete_Data_3_1035;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        713: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        714: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        715: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        716: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        717: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        718: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        719: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        720: begin
          delete_root_1080 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        721: begin
          delete_freeNext_9_index_196 <= delete_root_1080;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        722: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        723: begin
          delete_next_1079 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_1080;
          delete_freeNext_10_value_198 <= delete_indexRight_1075;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_1081 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        724: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_1075;
          delete_stuckIsFree_11_value_200 <= delete_isFree_1081;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        725: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        726: begin
          delete_freeNext_10_index_197 <= delete_indexRight_1075;
          delete_freeNext_10_value_198 <= delete_next_1079;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        727: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        728: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        729: begin
          delete_pc <= 730;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2490:Else|  Chip.java:0620:<init>|  Btree.java:2465:<init>|  Btree.java:2464:Then|  Chip.java:0610:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        730: begin
          delete_pc <= 829;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        731: begin
          if (delete_size_76 == 0) begin
            delete_pc <= 829;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        732: begin
          delete_index1_104 <= delete_size_76;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2497:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        733: begin
          delete_index1_104 <= delete_index1_104-1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0813:<init>|  Chip.java:0812:Dec|  Btree.java:2498:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        734: begin
          if (delete_index1_104 == 0) begin
            delete_pc <= 828;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        735: begin
          delete_index1_104 <= delete_index1_104-1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0813:<init>|  Chip.java:0812:Dec|  Btree.java:2505:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        736: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 780;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        737: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_1138 <= delete_Data_0_82;
              delete_indexRight_1139 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_1138 <= delete_Data_1_86;
              delete_indexRight_1139 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_1138 <= delete_Data_2_90;
              delete_indexRight_1139 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        738: begin
          delete_index_1082 <= delete_indexLeft_1138;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        739: begin
          delete_stuckSize_5_index_32 <= delete_index_1082;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_1082;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_1082;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_1082;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        740: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        741: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        742: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        743: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        744: begin
          delete_size_1083 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_1084 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_1086 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_1089 <= stuckData_stuckData_3_result_0;
          delete_Key_1_1090 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_1093 <= stuckData_stuckData_3_result_1;
          delete_Key_2_1094 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_1097 <= stuckData_stuckData_3_result_2;
          delete_Key_3_1098 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_1101 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        745: begin
          delete_index_1109 <= delete_indexRight_1139;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        746: begin
          delete_stuckSize_5_index_32 <= delete_index_1109;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_1109;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_1109;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_1109;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        747: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        748: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        749: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        750: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        751: begin
          delete_size_1110 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_1111 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_1113 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_1116 <= stuckData_stuckData_3_result_0;
          delete_Key_1_1117 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_1120 <= stuckData_stuckData_3_result_1;
          delete_Key_2_1121 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_1124 <= stuckData_stuckData_3_result_2;
          delete_Key_3_1125 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_1128 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        752: begin
          if (delete_isLeaf_1084 == 0) begin
            delete_pc <= 780;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        753: begin
          if (delete_isLeaf_1111 == 0) begin
            delete_pc <= 779;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        754: begin
          delete_MergeSuccess_1108 <= 0;
          case (delete_size_1083)
            0: begin
              case (delete_size_1110)
                0: begin
                  delete_size_1083 <= delete_size_1083 + 0;
                  delete_MergeSuccess_1108 <= 1;
                end
                1: begin
                  delete_Key_0_1086 <= delete_Key_0_1113;
                  delete_Data_0_1089 <= delete_Data_0_1116;
                  delete_size_1083 <= delete_size_1083 + 1;
                  delete_MergeSuccess_1108 <= 1;
                end
                2: begin
                  delete_Key_0_1086 <= delete_Key_0_1113;
                  delete_Data_0_1089 <= delete_Data_0_1116;
                  delete_Key_1_1090 <= delete_Key_1_1117;
                  delete_Data_1_1093 <= delete_Data_1_1120;
                  delete_size_1083 <= delete_size_1083 + 2;
                  delete_MergeSuccess_1108 <= 1;
                end
                3: begin
                  delete_Key_0_1086 <= delete_Key_0_1113;
                  delete_Data_0_1089 <= delete_Data_0_1116;
                  delete_Key_1_1090 <= delete_Key_1_1117;
                  delete_Data_1_1093 <= delete_Data_1_1120;
                  delete_Key_2_1094 <= delete_Key_2_1121;
                  delete_Data_2_1097 <= delete_Data_2_1124;
                  delete_size_1083 <= delete_size_1083 + 3;
                  delete_MergeSuccess_1108 <= 1;
                end
                4: begin
                  delete_Key_0_1086 <= delete_Key_0_1113;
                  delete_Data_0_1089 <= delete_Data_0_1116;
                  delete_Key_1_1090 <= delete_Key_1_1117;
                  delete_Data_1_1093 <= delete_Data_1_1120;
                  delete_Key_2_1094 <= delete_Key_2_1121;
                  delete_Data_2_1097 <= delete_Data_2_1124;
                  delete_Key_3_1098 <= delete_Key_3_1125;
                  delete_Data_3_1101 <= delete_Data_3_1128;
                  delete_size_1083 <= delete_size_1083 + 4;
                  delete_MergeSuccess_1108 <= 1;
                end
              endcase
            end
            1: begin
              case (delete_size_1110)
                0: begin
                  delete_size_1083 <= delete_size_1083 + 0;
                  delete_MergeSuccess_1108 <= 1;
                end
                1: begin
                  delete_Key_1_1090 <= delete_Key_0_1113;
                  delete_Data_1_1093 <= delete_Data_0_1116;
                  delete_size_1083 <= delete_size_1083 + 1;
                  delete_MergeSuccess_1108 <= 1;
                end
                2: begin
                  delete_Key_1_1090 <= delete_Key_0_1113;
                  delete_Data_1_1093 <= delete_Data_0_1116;
                  delete_Key_2_1094 <= delete_Key_1_1117;
                  delete_Data_2_1097 <= delete_Data_1_1120;
                  delete_size_1083 <= delete_size_1083 + 2;
                  delete_MergeSuccess_1108 <= 1;
                end
                3: begin
                  delete_Key_1_1090 <= delete_Key_0_1113;
                  delete_Data_1_1093 <= delete_Data_0_1116;
                  delete_Key_2_1094 <= delete_Key_1_1117;
                  delete_Data_2_1097 <= delete_Data_1_1120;
                  delete_Key_3_1098 <= delete_Key_2_1121;
                  delete_Data_3_1101 <= delete_Data_2_1124;
                  delete_size_1083 <= delete_size_1083 + 3;
                  delete_MergeSuccess_1108 <= 1;
                end
              endcase
            end
            2: begin
              case (delete_size_1110)
                0: begin
                  delete_size_1083 <= delete_size_1083 + 0;
                  delete_MergeSuccess_1108 <= 1;
                end
                1: begin
                  delete_Key_2_1094 <= delete_Key_0_1113;
                  delete_Data_2_1097 <= delete_Data_0_1116;
                  delete_size_1083 <= delete_size_1083 + 1;
                  delete_MergeSuccess_1108 <= 1;
                end
                2: begin
                  delete_Key_2_1094 <= delete_Key_0_1113;
                  delete_Data_2_1097 <= delete_Data_0_1116;
                  delete_Key_3_1098 <= delete_Key_1_1117;
                  delete_Data_3_1101 <= delete_Data_1_1120;
                  delete_size_1083 <= delete_size_1083 + 2;
                  delete_MergeSuccess_1108 <= 1;
                end
              endcase
            end
            3: begin
              case (delete_size_1110)
                0: begin
                  delete_size_1083 <= delete_size_1083 + 0;
                  delete_MergeSuccess_1108 <= 1;
                end
                1: begin
                  delete_Key_3_1098 <= delete_Key_0_1113;
                  delete_Data_3_1101 <= delete_Data_0_1116;
                  delete_size_1083 <= delete_size_1083 + 1;
                  delete_MergeSuccess_1108 <= 1;
                end
              endcase
            end
            4: begin
              case (delete_size_1110)
                0: begin
                  delete_size_1083 <= delete_size_1083 + 0;
                  delete_MergeSuccess_1108 <= 1;
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        755: begin
          if (delete_MergeSuccess_1108 == 0) begin
            delete_pc <= 778;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        756: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        757: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        758: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_1138;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_1138;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_1138;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_1138;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        759: begin
          delete_success_1141 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        760: begin
          delete_stuckSize_6_index_33 <= delete_index_1082;
          delete_stuckSize_6_value_34 <= delete_size_1083;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_1082;
          delete_stuckKeys_2_value_22 <= delete_Key_0_1086;
          delete_stuckKeys_2_value_23 <= delete_Key_1_1090;
          delete_stuckKeys_2_value_24 <= delete_Key_2_1094;
          delete_stuckKeys_2_value_25 <= delete_Key_3_1098;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_1082;
          delete_stuckData_4_value_28 <= delete_Data_0_1089;
          delete_stuckData_4_value_29 <= delete_Data_1_1093;
          delete_stuckData_4_value_30 <= delete_Data_2_1097;
          delete_stuckData_4_value_31 <= delete_Data_3_1101;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        761: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        762: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        763: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        764: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        765: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        766: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        767: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        768: begin
          delete_root_1144 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        769: begin
          delete_freeNext_9_index_196 <= delete_root_1144;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        770: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        771: begin
          delete_next_1143 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_1144;
          delete_freeNext_10_value_198 <= delete_indexRight_1139;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_1145 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        772: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_1139;
          delete_stuckIsFree_11_value_200 <= delete_isFree_1145;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        773: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        774: begin
          delete_freeNext_10_index_197 <= delete_indexRight_1139;
          delete_freeNext_10_value_198 <= delete_next_1143;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        775: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        776: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        777: begin
          delete_pc <= 778;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        778: begin
          delete_pc <= 779;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        779: begin
          delete_pc <= 780;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2506:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        780: begin
          if (delete_position_102 == 0 && delete_size_76 > 1) begin
            delete_pc <= delete_pc + 1;
          end
          else begin
            if (delete_position_102 == 0 || delete_size_76 < 1) begin
              delete_pc <= 827;
            end
            else begin
              delete_pc <= delete_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        781: begin
          delete_success_1207 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        782: begin
          case (delete_index1_104)
            0: begin
              delete_indexLeft_1204 <= delete_Data_0_82;
              delete_indexRight_1205 <= delete_Data_1_86;
            end
            1: begin
              delete_indexLeft_1204 <= delete_Data_1_86;
              delete_indexRight_1205 <= delete_Data_2_90;
            end
            2: begin
              delete_indexLeft_1204 <= delete_Data_2_90;
              delete_indexRight_1205 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        783: begin
          delete_index_1146 <= delete_indexLeft_1204;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        784: begin
          delete_stuckSize_5_index_32 <= delete_index_1146;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_1146;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_1146;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_1146;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        785: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        786: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        787: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        788: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        789: begin
          delete_size_1147 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_1148 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_1150 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_1153 <= stuckData_stuckData_3_result_0;
          delete_Key_1_1154 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_1157 <= stuckData_stuckData_3_result_1;
          delete_Key_2_1158 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_1161 <= stuckData_stuckData_3_result_2;
          delete_Key_3_1162 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_1165 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        790: begin
          delete_index_1173 <= delete_indexRight_1205;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        791: begin
          delete_stuckSize_5_index_32 <= delete_index_1173;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_1173;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_1173;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_1173;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        792: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        793: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        794: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        795: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        796: begin
          delete_size_1174 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_1175 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_1177 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_1180 <= stuckData_stuckData_3_result_0;
          delete_Key_1_1181 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_1184 <= stuckData_stuckData_3_result_1;
          delete_Key_2_1185 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_1188 <= stuckData_stuckData_3_result_2;
          delete_Key_3_1189 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_1192 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        797: begin
          if (delete_isLeaf_1148 == 0) begin
            delete_pc <= 799;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        798: begin
          delete_pc <= 827;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        799: begin
          if (delete_isLeaf_1175 == 0) begin
            delete_pc <= 801;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        800: begin
          delete_pc <= 827;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        801: begin
          case (delete_index1_104)
            0: begin
              delete_midKey_1206 <= delete_Key_0_79;
            end
            1: begin
              delete_midKey_1206 <= delete_Key_1_83;
            end
            2: begin
              delete_midKey_1206 <= delete_Key_2_87;
            end
            3: begin
              delete_midKey_1206 <= delete_Key_3_91;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        802: begin
          delete_MergeSuccess_1172 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        803: begin
          case (delete_size_1147)
            0: begin
              case (delete_size_1174)
                0: begin
                  delete_Key_0_1150 <= delete_midKey_1206;
                  delete_Data_1_1157 <= delete_Data_0_1180;
                  delete_size_1147 <= delete_size_1147 + 1;
                  delete_MergeSuccess_1172 <= 1;
                end
                1: begin
                  delete_Key_0_1150 <= delete_midKey_1206;
                  delete_Key_1_1154 <= delete_Key_0_1177;
                  delete_Data_1_1157 <= delete_Data_0_1180;
                  delete_Data_2_1161 <= delete_Data_1_1184;
                  delete_size_1147 <= delete_size_1147 + 2;
                  delete_MergeSuccess_1172 <= 1;
                end
                2: begin
                  delete_Key_0_1150 <= delete_midKey_1206;
                  delete_Key_1_1154 <= delete_Key_0_1177;
                  delete_Data_1_1157 <= delete_Data_0_1180;
                  delete_Key_2_1158 <= delete_Key_1_1181;
                  delete_Data_2_1161 <= delete_Data_1_1184;
                  delete_Data_3_1165 <= delete_Data_2_1188;
                  delete_size_1147 <= delete_size_1147 + 3;
                  delete_MergeSuccess_1172 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (delete_size_1174)
                0: begin
                  delete_Key_1_1154 <= delete_midKey_1206;
                  delete_Data_2_1161 <= delete_Data_0_1180;
                  delete_size_1147 <= delete_size_1147 + 1;
                  delete_MergeSuccess_1172 <= 1;
                end
                1: begin
                  delete_Key_1_1154 <= delete_midKey_1206;
                  delete_Key_2_1158 <= delete_Key_0_1177;
                  delete_Data_2_1161 <= delete_Data_0_1180;
                  delete_Data_3_1165 <= delete_Data_1_1184;
                  delete_size_1147 <= delete_size_1147 + 2;
                  delete_MergeSuccess_1172 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (delete_size_1174)
                0: begin
                  delete_Key_2_1158 <= delete_midKey_1206;
                  delete_Data_3_1165 <= delete_Data_0_1180;
                  delete_size_1147 <= delete_size_1147 + 1;
                  delete_MergeSuccess_1172 <= 1;
                end
                1: begin
                end
                2: begin
                end
              endcase
            end
            3: begin
              case (delete_size_1174)
                0: begin
                end
                1: begin
                end
              endcase
            end
            4: begin
              case (delete_size_1174)
                0: begin
                end
              endcase
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        804: begin
          if (delete_MergeSuccess_1172 == 0) begin
            delete_pc <= 827;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        805: begin
          delete_size_76 <= delete_size_76-1;
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          if (0>= delete_index1_104) begin
            delete_Key_0_79 <= delete_Key_1_83;
            delete_Data_0_82 <= delete_Data_1_86;
          end
          if (1>= delete_index1_104) begin
            delete_Key_1_83 <= delete_Key_2_87;
            delete_Data_1_86 <= delete_Data_2_90;
          end
          if (2>= delete_index1_104) begin
            delete_Key_2_87 <= delete_Key_3_91;
            delete_Data_2_90 <= delete_Data_3_94;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        806: begin
          case (delete_index1_104)
            0: begin
              delete_Key_96 <= delete_Key_0_79;
              delete_Data_98 <= delete_Data_0_82;
            end
            1: begin
              delete_Key_96 <= delete_Key_1_83;
              delete_Data_98 <= delete_Data_1_86;
            end
            2: begin
              delete_Key_96 <= delete_Key_2_87;
              delete_Data_98 <= delete_Data_2_90;
            end
            3: begin
              delete_Key_96 <= delete_Key_3_91;
              delete_Data_98 <= delete_Data_3_94;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        807: begin
          if (delete_index1_104 == delete_size_76) begin
            delete_size_76 <= delete_size_76+1;
          end
          case (delete_index1_104)
            0: begin
              delete_Key_0_79 <= delete_Key_96;
              delete_Data_0_82 <= delete_indexLeft_1204;
            end
            1: begin
              delete_Key_1_83 <= delete_Key_96;
              delete_Data_1_86 <= delete_indexLeft_1204;
            end
            2: begin
              delete_Key_2_87 <= delete_Key_96;
              delete_Data_2_90 <= delete_indexLeft_1204;
            end
            3: begin
              delete_Key_3_91 <= delete_Key_96;
              delete_Data_3_94 <= delete_indexLeft_1204;
            end
          endcase
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        808: begin
          delete_success_1207 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        809: begin
          delete_stuckSize_6_index_33 <= delete_index_1146;
          delete_stuckSize_6_value_34 <= delete_size_1147;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_1146;
          delete_stuckKeys_2_value_22 <= delete_Key_0_1150;
          delete_stuckKeys_2_value_23 <= delete_Key_1_1154;
          delete_stuckKeys_2_value_24 <= delete_Key_2_1158;
          delete_stuckKeys_2_value_25 <= delete_Key_3_1162;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_1146;
          delete_stuckData_4_value_28 <= delete_Data_0_1153;
          delete_stuckData_4_value_29 <= delete_Data_1_1157;
          delete_stuckData_4_value_30 <= delete_Data_2_1161;
          delete_stuckData_4_value_31 <= delete_Data_3_1165;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        810: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        811: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        812: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        813: begin
          delete_stuckSize_6_index_33 <= delete_index_75;
          delete_stuckSize_6_value_34 <= delete_size_76;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          delete_stuckKeys_2_index_21 <= delete_index_75;
          delete_stuckKeys_2_value_22 <= delete_Key_0_79;
          delete_stuckKeys_2_value_23 <= delete_Key_1_83;
          delete_stuckKeys_2_value_24 <= delete_Key_2_87;
          delete_stuckKeys_2_value_25 <= delete_Key_3_91;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          delete_stuckData_4_index_27 <= delete_index_75;
          delete_stuckData_4_value_28 <= delete_Data_0_82;
          delete_stuckData_4_value_29 <= delete_Data_1_86;
          delete_stuckData_4_value_30 <= delete_Data_2_90;
          delete_stuckData_4_value_31 <= delete_Data_3_94;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        814: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        815: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        816: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        817: begin
          delete_root_1210 <= 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        818: begin
          delete_freeNext_9_index_196 <= delete_root_1210;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        819: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        820: begin
          delete_next_1209 <= freeNext_freeNext_9_result_0;
          delete_freeNext_10_index_197 <= delete_root_1210;
          delete_freeNext_10_value_198 <= delete_indexRight_1205;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_isFree_1211 <= 1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        821: begin
          delete_stuckIsFree_11_index_199 <= delete_indexRight_1205;
          delete_stuckIsFree_11_value_200 <= delete_isFree_1211;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        822: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        823: begin
          delete_freeNext_10_index_197 <= delete_indexRight_1205;
          delete_freeNext_10_value_198 <= delete_next_1209;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        824: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        825: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        826: begin
          delete_pc <= 827;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2507:Then|  Chip.java:0610:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        827: begin
          delete_pc <= 828;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2504:<init>|  Btree.java:2503:Then|  Chip.java:0610:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        828: begin
          delete_pc <= 829;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2496:<init>|  Btree.java:2495:Else|  Chip.java:0620:<init>|  Btree.java:2463:<init>|  Btree.java:2462:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        829: begin
          delete_index_75 <= delete_position_102;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        830: begin
          delete_stuckSize_5_index_32 <= delete_index_75;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_75;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_75;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_75;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        831: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        832: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        833: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        834: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        835: begin
          delete_size_76 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_77 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_79 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_82 <= stuckData_stuckData_3_result_0;
          delete_Key_1_83 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_86 <= stuckData_stuckData_3_result_1;
          delete_Key_2_87 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_90 <= stuckData_stuckData_3_result_2;
          delete_Key_3_91 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_94 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2515:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        836: begin
          delete_KeyCompares_0_80 <= delete_k_46 <= delete_Key_0_79 && 0 < delete_size_76;
          delete_KeyCollapse_0_81 <= 0;
          delete_KeyCompares_1_84 <= delete_k_46 >  delete_Key_0_79 && delete_k_46 <= delete_Key_1_83 && 1 < delete_size_76;
          delete_KeyCollapse_1_85 <= 1;
          delete_KeyCompares_2_88 <= delete_k_46 >  delete_Key_1_83 && delete_k_46 <= delete_Key_2_87 && 2 < delete_size_76;
          delete_KeyCollapse_2_89 <= 2;
          delete_KeyCompares_3_92 <= delete_k_46 >  delete_Key_2_87 && delete_k_46 <= delete_Key_3_91 && 3 < delete_size_76;
          delete_KeyCollapse_3_93 <= 3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2516:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        837: begin
          if (delete_KeyCompares_1_84) begin
            delete_KeyCompares_0_80 <= 1;
            delete_KeyCollapse_0_81 <= delete_KeyCollapse_1_85;
          end
          if (delete_KeyCompares_3_92) begin
            delete_KeyCompares_2_88 <= 1;
            delete_KeyCollapse_2_89 <= delete_KeyCollapse_3_93;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2516:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        838: begin
          if (delete_KeyCompares_2_88) begin
            delete_KeyCompares_0_80 <= 1;
            delete_KeyCollapse_0_81 <= delete_KeyCollapse_2_89;
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2516:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        839: begin
          if (delete_KeyCompares_0_80) begin
            delete_Found_95 <= 1;
            case (delete_KeyCollapse_0_81)
              0: begin
                delete_StuckIndex_100 <= 0;
                delete_FoundKey_97 <= delete_Key_0_79;
                delete_Data_98 <= delete_Data_0_82;
              end
              1: begin
                delete_StuckIndex_100 <= 1;
                delete_FoundKey_97 <= delete_Key_1_83;
                delete_Data_98 <= delete_Data_1_86;
              end
              2: begin
                delete_StuckIndex_100 <= 2;
                delete_FoundKey_97 <= delete_Key_2_87;
                delete_Data_98 <= delete_Data_2_90;
              end
              3: begin
                delete_StuckIndex_100 <= 3;
                delete_FoundKey_97 <= delete_Key_3_91;
                delete_Data_98 <= delete_Data_3_94;
              end
            endcase
          end
          else begin
            delete_Found_95 <= 0;
            case (delete_size_76)
              0: begin
                delete_StuckIndex_100 <= 0;
                delete_Data_98 <= delete_Data_0_82;
              end
              1: begin
                delete_StuckIndex_100 <= 1;
                delete_Data_98 <= delete_Data_1_86;
              end
              2: begin
                delete_StuckIndex_100 <= 2;
                delete_Data_98 <= delete_Data_2_90;
              end
              3: begin
                delete_StuckIndex_100 <= 3;
                delete_Data_98 <= delete_Data_3_94;
              end
            endcase
          end
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2516:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        840: begin
          delete_position_102 <= delete_Data_98;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2517:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        841: begin
          delete_index_75 <= delete_position_102;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        842: begin
          delete_stuckSize_5_index_32 <= delete_index_75;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          delete_stuckIsLeaf_7_index_35 <= delete_index_75;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          delete_stuckKeys_1_index_20 <= delete_index_75;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          delete_stuckData_3_index_26 <= delete_index_75;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        843: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        844: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        845: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        846: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        847: begin
          delete_size_76 <= stuckSize_stuckSize_5_result_0;
          delete_isLeaf_77 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          delete_Key_0_79 <= stuckKeys_stuckKeys_1_result_0;
          delete_Data_0_82 <= stuckData_stuckData_3_result_0;
          delete_Key_1_83 <= stuckKeys_stuckKeys_1_result_1;
          delete_Data_1_86 <= stuckData_stuckData_3_result_1;
          delete_Key_2_87 <= stuckKeys_stuckKeys_1_result_2;
          delete_Data_2_90 <= stuckData_stuckData_3_result_2;
          delete_Key_3_91 <= stuckKeys_stuckKeys_1_result_3;
          delete_Data_3_94 <= stuckData_stuckData_3_result_3;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2519:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        848: begin
          if (delete_isLeaf_77 == 0) begin
            delete_pc <= 851;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2522:<init>|  Btree.java:2521:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        849: begin
          delete_pc <= 852;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2523:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2522:<init>|  Btree.java:2521:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        850: begin
          delete_pc <= 852;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2522:<init>|  Btree.java:2521:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        851: begin
          delete_pc <= 166;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2526:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2522:<init>|  Btree.java:2521:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2634:Then|  Chip.java:0610:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        852: begin
          delete_pc <= 853;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2624:<init>|  Btree.java:2623:code|  Chip.java:0530:<init>|  Btree.java:2621:<init>|  Btree.java:2620:delete|  Btree.java:5325:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        853: begin
          delete_l_47 <= delete_i_45< 32 ? 1 : 0;
          delete_pc <= delete_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:5327:<init>|  Btree.java:5326:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        854: begin
          if (delete_l_47 >  0) begin
            delete_pc <= 1;
          end
          else begin
            delete_pc <= delete_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0578:<init>|  Chip.java:0577:GONotZero|  Btree.java:5335:code|  Chip.java:0530:<init>|  Btree.java:5309:<init>|  Btree.java:5308:test_delete_descending|  Btree.java:6876:newTests|  Btree.java:6882:main|");
            $fclose(f);
          end
        end
        default: delete_stop <= 1;
      endcase
    end
  end
  task chipPrint;
    begin
      integer o;
      o = $fopen("verilog/trace_verilog.txt", "a");
      if (!o) o = $fopen("../verilog/trace_verilog.txt", "a");
      if (!o) $display("Cannot create trace folder: verilog/trace_verilog.txt");
      $fwrite(o, "Chip: %-16s step: %1d, maxSteps: %1d, running: %1d\n", "Btree", step, maxSteps, !stop);
      $fwrite(o, "  Processes:\n");

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 0, "stuckIsLeaf", 1, stuckIsLeaf_pc, stuckIsLeaf_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsLeaf_memory[0]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[1]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[2]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[3]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[4]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[5]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[6]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[7]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[8]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[9]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[10]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[11]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[12]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[13]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[14]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[15]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[16]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[17]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[18]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[19]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[20]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[21]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[22]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[23]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[24]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[25]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[26]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[27]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[28]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[29]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[30]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckIsLeaf_7", stuckIsLeaf_7_requestedAt, stuckIsLeaf_7_finishedAt, stuckIsLeaf_stuckIsLeaf_7_returnCode, (stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step), (stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckIsLeaf_7_index_35", delete_stuckIsLeaf_7_index_35);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsLeaf_8", stuckIsLeaf_8_requestedAt, stuckIsLeaf_8_finishedAt, stuckIsLeaf_stuckIsLeaf_8_returnCode, (stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step), (stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckIsLeaf_8_index_36", delete_stuckIsLeaf_8_index_36);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckIsLeaf_8_value_37", delete_stuckIsLeaf_8_value_37);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 1, "stuckIsFree", 1, stuckIsFree_pc, stuckIsFree_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsFree_memory[0]);
      $fwrite(o, ", %2d", stuckIsFree_memory[1]);
      $fwrite(o, ", %2d", stuckIsFree_memory[2]);
      $fwrite(o, ", %2d", stuckIsFree_memory[3]);
      $fwrite(o, ", %2d", stuckIsFree_memory[4]);
      $fwrite(o, ", %2d", stuckIsFree_memory[5]);
      $fwrite(o, ", %2d", stuckIsFree_memory[6]);
      $fwrite(o, ", %2d", stuckIsFree_memory[7]);
      $fwrite(o, ", %2d", stuckIsFree_memory[8]);
      $fwrite(o, ", %2d", stuckIsFree_memory[9]);
      $fwrite(o, ", %2d", stuckIsFree_memory[10]);
      $fwrite(o, ", %2d", stuckIsFree_memory[11]);
      $fwrite(o, ", %2d", stuckIsFree_memory[12]);
      $fwrite(o, ", %2d", stuckIsFree_memory[13]);
      $fwrite(o, ", %2d", stuckIsFree_memory[14]);
      $fwrite(o, ", %2d", stuckIsFree_memory[15]);
      $fwrite(o, ", %2d", stuckIsFree_memory[16]);
      $fwrite(o, ", %2d", stuckIsFree_memory[17]);
      $fwrite(o, ", %2d", stuckIsFree_memory[18]);
      $fwrite(o, ", %2d", stuckIsFree_memory[19]);
      $fwrite(o, ", %2d", stuckIsFree_memory[20]);
      $fwrite(o, ", %2d", stuckIsFree_memory[21]);
      $fwrite(o, ", %2d", stuckIsFree_memory[22]);
      $fwrite(o, ", %2d", stuckIsFree_memory[23]);
      $fwrite(o, ", %2d", stuckIsFree_memory[24]);
      $fwrite(o, ", %2d", stuckIsFree_memory[25]);
      $fwrite(o, ", %2d", stuckIsFree_memory[26]);
      $fwrite(o, ", %2d", stuckIsFree_memory[27]);
      $fwrite(o, ", %2d", stuckIsFree_memory[28]);
      $fwrite(o, ", %2d", stuckIsFree_memory[29]);
      $fwrite(o, ", %2d", stuckIsFree_memory[30]);
      $fwrite(o, ", %2d", stuckIsFree_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsFree_11", stuckIsFree_11_requestedAt, stuckIsFree_11_finishedAt, stuckIsFree_stuckIsFree_11_returnCode, (stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step), (stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckIsFree_11_index_199", delete_stuckIsFree_11_index_199);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckIsFree_11_value_200", delete_stuckIsFree_11_value_200);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 2, "freeNext", 1, freeNext_pc, freeNext_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 6, 1);
      $fwrite(o, "        %2d", freeNext_memory[0]);
      $fwrite(o, ", %2d", freeNext_memory[1]);
      $fwrite(o, ", %2d", freeNext_memory[2]);
      $fwrite(o, ", %2d", freeNext_memory[3]);
      $fwrite(o, ", %2d", freeNext_memory[4]);
      $fwrite(o, ", %2d", freeNext_memory[5]);
      $fwrite(o, ", %2d", freeNext_memory[6]);
      $fwrite(o, ", %2d", freeNext_memory[7]);
      $fwrite(o, ", %2d", freeNext_memory[8]);
      $fwrite(o, ", %2d", freeNext_memory[9]);
      $fwrite(o, ", %2d", freeNext_memory[10]);
      $fwrite(o, ", %2d", freeNext_memory[11]);
      $fwrite(o, ", %2d", freeNext_memory[12]);
      $fwrite(o, ", %2d", freeNext_memory[13]);
      $fwrite(o, ", %2d", freeNext_memory[14]);
      $fwrite(o, ", %2d", freeNext_memory[15]);
      $fwrite(o, ", %2d", freeNext_memory[16]);
      $fwrite(o, ", %2d", freeNext_memory[17]);
      $fwrite(o, ", %2d", freeNext_memory[18]);
      $fwrite(o, ", %2d", freeNext_memory[19]);
      $fwrite(o, ", %2d", freeNext_memory[20]);
      $fwrite(o, ", %2d", freeNext_memory[21]);
      $fwrite(o, ", %2d", freeNext_memory[22]);
      $fwrite(o, ", %2d", freeNext_memory[23]);
      $fwrite(o, ", %2d", freeNext_memory[24]);
      $fwrite(o, ", %2d", freeNext_memory[25]);
      $fwrite(o, ", %2d", freeNext_memory[26]);
      $fwrite(o, ", %2d", freeNext_memory[27]);
      $fwrite(o, ", %2d", freeNext_memory[28]);
      $fwrite(o, ", %2d", freeNext_memory[29]);
      $fwrite(o, ", %2d", freeNext_memory[30]);
      $fwrite(o, ", %2d", freeNext_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "freeNext_9", freeNext_9_requestedAt, freeNext_9_finishedAt, freeNext_freeNext_9_returnCode, (freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step), (freeNext_9_requestedAt < freeNext_9_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_freeNext_9_index_196", delete_freeNext_9_index_196);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "freeNext_10", freeNext_10_requestedAt, freeNext_10_finishedAt, freeNext_freeNext_10_returnCode, (freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step), (freeNext_10_requestedAt < freeNext_10_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_freeNext_10_index_197", delete_freeNext_10_index_197);

      $fwrite(o, "            %-38s = %1d\n", "delete_freeNext_10_value_198", delete_freeNext_10_value_198);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 3, "stuckSize", 1, stuckSize_pc, stuckSize_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 3, 1);
      $fwrite(o, "        %2d", stuckSize_memory[0]);
      $fwrite(o, ", %2d", stuckSize_memory[1]);
      $fwrite(o, ", %2d", stuckSize_memory[2]);
      $fwrite(o, ", %2d", stuckSize_memory[3]);
      $fwrite(o, ", %2d", stuckSize_memory[4]);
      $fwrite(o, ", %2d", stuckSize_memory[5]);
      $fwrite(o, ", %2d", stuckSize_memory[6]);
      $fwrite(o, ", %2d", stuckSize_memory[7]);
      $fwrite(o, ", %2d", stuckSize_memory[8]);
      $fwrite(o, ", %2d", stuckSize_memory[9]);
      $fwrite(o, ", %2d", stuckSize_memory[10]);
      $fwrite(o, ", %2d", stuckSize_memory[11]);
      $fwrite(o, ", %2d", stuckSize_memory[12]);
      $fwrite(o, ", %2d", stuckSize_memory[13]);
      $fwrite(o, ", %2d", stuckSize_memory[14]);
      $fwrite(o, ", %2d", stuckSize_memory[15]);
      $fwrite(o, ", %2d", stuckSize_memory[16]);
      $fwrite(o, ", %2d", stuckSize_memory[17]);
      $fwrite(o, ", %2d", stuckSize_memory[18]);
      $fwrite(o, ", %2d", stuckSize_memory[19]);
      $fwrite(o, ", %2d", stuckSize_memory[20]);
      $fwrite(o, ", %2d", stuckSize_memory[21]);
      $fwrite(o, ", %2d", stuckSize_memory[22]);
      $fwrite(o, ", %2d", stuckSize_memory[23]);
      $fwrite(o, ", %2d", stuckSize_memory[24]);
      $fwrite(o, ", %2d", stuckSize_memory[25]);
      $fwrite(o, ", %2d", stuckSize_memory[26]);
      $fwrite(o, ", %2d", stuckSize_memory[27]);
      $fwrite(o, ", %2d", stuckSize_memory[28]);
      $fwrite(o, ", %2d", stuckSize_memory[29]);
      $fwrite(o, ", %2d", stuckSize_memory[30]);
      $fwrite(o, ", %2d", stuckSize_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckSize_5", stuckSize_5_requestedAt, stuckSize_5_finishedAt, stuckSize_stuckSize_5_returnCode, (stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step), (stuckSize_5_requestedAt < stuckSize_5_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckSize_5_index_32", delete_stuckSize_5_index_32);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckSize_6", stuckSize_6_requestedAt, stuckSize_6_finishedAt, stuckSize_stuckSize_6_returnCode, (stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step), (stuckSize_6_requestedAt < stuckSize_6_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckSize_6_index_33", delete_stuckSize_6_index_33);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckSize_6_value_34", delete_stuckSize_6_value_34);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 4, "stuckKeys", 1, stuckKeys_pc, stuckKeys_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckKeys_memory[0]);
      $fwrite(o, ", %2d", stuckKeys_memory[1]);
      $fwrite(o, ", %2d", stuckKeys_memory[2]);
      $fwrite(o, ", %2d", stuckKeys_memory[3]);
      $fwrite(o, ", %2d", stuckKeys_memory[4]);
      $fwrite(o, ", %2d", stuckKeys_memory[5]);
      $fwrite(o, ", %2d", stuckKeys_memory[6]);
      $fwrite(o, ", %2d", stuckKeys_memory[7]);
      $fwrite(o, ", %2d", stuckKeys_memory[8]);
      $fwrite(o, ", %2d", stuckKeys_memory[9]);
      $fwrite(o, ", %2d", stuckKeys_memory[10]);
      $fwrite(o, ", %2d", stuckKeys_memory[11]);
      $fwrite(o, ", %2d", stuckKeys_memory[12]);
      $fwrite(o, ", %2d", stuckKeys_memory[13]);
      $fwrite(o, ", %2d", stuckKeys_memory[14]);
      $fwrite(o, ", %2d", stuckKeys_memory[15]);
      $fwrite(o, ", %2d", stuckKeys_memory[16]);
      $fwrite(o, ", %2d", stuckKeys_memory[17]);
      $fwrite(o, ", %2d", stuckKeys_memory[18]);
      $fwrite(o, ", %2d", stuckKeys_memory[19]);
      $fwrite(o, ", %2d", stuckKeys_memory[20]);
      $fwrite(o, ", %2d", stuckKeys_memory[21]);
      $fwrite(o, ", %2d", stuckKeys_memory[22]);
      $fwrite(o, ", %2d", stuckKeys_memory[23]);
      $fwrite(o, ", %2d", stuckKeys_memory[24]);
      $fwrite(o, ", %2d", stuckKeys_memory[25]);
      $fwrite(o, ", %2d", stuckKeys_memory[26]);
      $fwrite(o, ", %2d", stuckKeys_memory[27]);
      $fwrite(o, ", %2d", stuckKeys_memory[28]);
      $fwrite(o, ", %2d", stuckKeys_memory[29]);
      $fwrite(o, ", %2d", stuckKeys_memory[30]);
      $fwrite(o, ", %2d", stuckKeys_memory[31]);
      $fwrite(o, ", %2d", stuckKeys_memory[32]);
      $fwrite(o, ", %2d", stuckKeys_memory[33]);
      $fwrite(o, ", %2d", stuckKeys_memory[34]);
      $fwrite(o, ", %2d", stuckKeys_memory[35]);
      $fwrite(o, ", %2d", stuckKeys_memory[36]);
      $fwrite(o, ", %2d", stuckKeys_memory[37]);
      $fwrite(o, ", %2d", stuckKeys_memory[38]);
      $fwrite(o, ", %2d", stuckKeys_memory[39]);
      $fwrite(o, ", %2d", stuckKeys_memory[40]);
      $fwrite(o, ", %2d", stuckKeys_memory[41]);
      $fwrite(o, ", %2d", stuckKeys_memory[42]);
      $fwrite(o, ", %2d", stuckKeys_memory[43]);
      $fwrite(o, ", %2d", stuckKeys_memory[44]);
      $fwrite(o, ", %2d", stuckKeys_memory[45]);
      $fwrite(o, ", %2d", stuckKeys_memory[46]);
      $fwrite(o, ", %2d", stuckKeys_memory[47]);
      $fwrite(o, ", %2d", stuckKeys_memory[48]);
      $fwrite(o, ", %2d", stuckKeys_memory[49]);
      $fwrite(o, ", %2d", stuckKeys_memory[50]);
      $fwrite(o, ", %2d", stuckKeys_memory[51]);
      $fwrite(o, ", %2d", stuckKeys_memory[52]);
      $fwrite(o, ", %2d", stuckKeys_memory[53]);
      $fwrite(o, ", %2d", stuckKeys_memory[54]);
      $fwrite(o, ", %2d", stuckKeys_memory[55]);
      $fwrite(o, ", %2d", stuckKeys_memory[56]);
      $fwrite(o, ", %2d", stuckKeys_memory[57]);
      $fwrite(o, ", %2d", stuckKeys_memory[58]);
      $fwrite(o, ", %2d", stuckKeys_memory[59]);
      $fwrite(o, ", %2d", stuckKeys_memory[60]);
      $fwrite(o, ", %2d", stuckKeys_memory[61]);
      $fwrite(o, ", %2d", stuckKeys_memory[62]);
      $fwrite(o, ", %2d", stuckKeys_memory[63]);
      $fwrite(o, ", %2d", stuckKeys_memory[64]);
      $fwrite(o, ", %2d", stuckKeys_memory[65]);
      $fwrite(o, ", %2d", stuckKeys_memory[66]);
      $fwrite(o, ", %2d", stuckKeys_memory[67]);
      $fwrite(o, ", %2d", stuckKeys_memory[68]);
      $fwrite(o, ", %2d", stuckKeys_memory[69]);
      $fwrite(o, ", %2d", stuckKeys_memory[70]);
      $fwrite(o, ", %2d", stuckKeys_memory[71]);
      $fwrite(o, ", %2d", stuckKeys_memory[72]);
      $fwrite(o, ", %2d", stuckKeys_memory[73]);
      $fwrite(o, ", %2d", stuckKeys_memory[74]);
      $fwrite(o, ", %2d", stuckKeys_memory[75]);
      $fwrite(o, ", %2d", stuckKeys_memory[76]);
      $fwrite(o, ", %2d", stuckKeys_memory[77]);
      $fwrite(o, ", %2d", stuckKeys_memory[78]);
      $fwrite(o, ", %2d", stuckKeys_memory[79]);
      $fwrite(o, ", %2d", stuckKeys_memory[80]);
      $fwrite(o, ", %2d", stuckKeys_memory[81]);
      $fwrite(o, ", %2d", stuckKeys_memory[82]);
      $fwrite(o, ", %2d", stuckKeys_memory[83]);
      $fwrite(o, ", %2d", stuckKeys_memory[84]);
      $fwrite(o, ", %2d", stuckKeys_memory[85]);
      $fwrite(o, ", %2d", stuckKeys_memory[86]);
      $fwrite(o, ", %2d", stuckKeys_memory[87]);
      $fwrite(o, ", %2d", stuckKeys_memory[88]);
      $fwrite(o, ", %2d", stuckKeys_memory[89]);
      $fwrite(o, ", %2d", stuckKeys_memory[90]);
      $fwrite(o, ", %2d", stuckKeys_memory[91]);
      $fwrite(o, ", %2d", stuckKeys_memory[92]);
      $fwrite(o, ", %2d", stuckKeys_memory[93]);
      $fwrite(o, ", %2d", stuckKeys_memory[94]);
      $fwrite(o, ", %2d", stuckKeys_memory[95]);
      $fwrite(o, ", %2d", stuckKeys_memory[96]);
      $fwrite(o, ", %2d", stuckKeys_memory[97]);
      $fwrite(o, ", %2d", stuckKeys_memory[98]);
      $fwrite(o, ", %2d", stuckKeys_memory[99]);
      $fwrite(o, ", %2d", stuckKeys_memory[100]);
      $fwrite(o, ", %2d", stuckKeys_memory[101]);
      $fwrite(o, ", %2d", stuckKeys_memory[102]);
      $fwrite(o, ", %2d", stuckKeys_memory[103]);
      $fwrite(o, ", %2d", stuckKeys_memory[104]);
      $fwrite(o, ", %2d", stuckKeys_memory[105]);
      $fwrite(o, ", %2d", stuckKeys_memory[106]);
      $fwrite(o, ", %2d", stuckKeys_memory[107]);
      $fwrite(o, ", %2d", stuckKeys_memory[108]);
      $fwrite(o, ", %2d", stuckKeys_memory[109]);
      $fwrite(o, ", %2d", stuckKeys_memory[110]);
      $fwrite(o, ", %2d", stuckKeys_memory[111]);
      $fwrite(o, ", %2d", stuckKeys_memory[112]);
      $fwrite(o, ", %2d", stuckKeys_memory[113]);
      $fwrite(o, ", %2d", stuckKeys_memory[114]);
      $fwrite(o, ", %2d", stuckKeys_memory[115]);
      $fwrite(o, ", %2d", stuckKeys_memory[116]);
      $fwrite(o, ", %2d", stuckKeys_memory[117]);
      $fwrite(o, ", %2d", stuckKeys_memory[118]);
      $fwrite(o, ", %2d", stuckKeys_memory[119]);
      $fwrite(o, ", %2d", stuckKeys_memory[120]);
      $fwrite(o, ", %2d", stuckKeys_memory[121]);
      $fwrite(o, ", %2d", stuckKeys_memory[122]);
      $fwrite(o, ", %2d", stuckKeys_memory[123]);
      $fwrite(o, ", %2d", stuckKeys_memory[124]);
      $fwrite(o, ", %2d", stuckKeys_memory[125]);
      $fwrite(o, ", %2d", stuckKeys_memory[126]);
      $fwrite(o, ", %2d", stuckKeys_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckKeys_1", stuckKeys_1_requestedAt, stuckKeys_1_finishedAt, stuckKeys_stuckKeys_1_returnCode, (stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step), (stuckKeys_1_requestedAt < stuckKeys_1_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckKeys_1_index_20", delete_stuckKeys_1_index_20);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckKeys_2", stuckKeys_2_requestedAt, stuckKeys_2_finishedAt, stuckKeys_stuckKeys_2_returnCode, (stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step), (stuckKeys_2_requestedAt < stuckKeys_2_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckKeys_2_index_21", delete_stuckKeys_2_index_21);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckKeys_2_value_22", delete_stuckKeys_2_value_22);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckKeys_2_value_23", delete_stuckKeys_2_value_23);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckKeys_2_value_24", delete_stuckKeys_2_value_24);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckKeys_2_value_25", delete_stuckKeys_2_value_25);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 5, "stuckData", 1, stuckData_pc, stuckData_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckData_memory[0]);
      $fwrite(o, ", %2d", stuckData_memory[1]);
      $fwrite(o, ", %2d", stuckData_memory[2]);
      $fwrite(o, ", %2d", stuckData_memory[3]);
      $fwrite(o, ", %2d", stuckData_memory[4]);
      $fwrite(o, ", %2d", stuckData_memory[5]);
      $fwrite(o, ", %2d", stuckData_memory[6]);
      $fwrite(o, ", %2d", stuckData_memory[7]);
      $fwrite(o, ", %2d", stuckData_memory[8]);
      $fwrite(o, ", %2d", stuckData_memory[9]);
      $fwrite(o, ", %2d", stuckData_memory[10]);
      $fwrite(o, ", %2d", stuckData_memory[11]);
      $fwrite(o, ", %2d", stuckData_memory[12]);
      $fwrite(o, ", %2d", stuckData_memory[13]);
      $fwrite(o, ", %2d", stuckData_memory[14]);
      $fwrite(o, ", %2d", stuckData_memory[15]);
      $fwrite(o, ", %2d", stuckData_memory[16]);
      $fwrite(o, ", %2d", stuckData_memory[17]);
      $fwrite(o, ", %2d", stuckData_memory[18]);
      $fwrite(o, ", %2d", stuckData_memory[19]);
      $fwrite(o, ", %2d", stuckData_memory[20]);
      $fwrite(o, ", %2d", stuckData_memory[21]);
      $fwrite(o, ", %2d", stuckData_memory[22]);
      $fwrite(o, ", %2d", stuckData_memory[23]);
      $fwrite(o, ", %2d", stuckData_memory[24]);
      $fwrite(o, ", %2d", stuckData_memory[25]);
      $fwrite(o, ", %2d", stuckData_memory[26]);
      $fwrite(o, ", %2d", stuckData_memory[27]);
      $fwrite(o, ", %2d", stuckData_memory[28]);
      $fwrite(o, ", %2d", stuckData_memory[29]);
      $fwrite(o, ", %2d", stuckData_memory[30]);
      $fwrite(o, ", %2d", stuckData_memory[31]);
      $fwrite(o, ", %2d", stuckData_memory[32]);
      $fwrite(o, ", %2d", stuckData_memory[33]);
      $fwrite(o, ", %2d", stuckData_memory[34]);
      $fwrite(o, ", %2d", stuckData_memory[35]);
      $fwrite(o, ", %2d", stuckData_memory[36]);
      $fwrite(o, ", %2d", stuckData_memory[37]);
      $fwrite(o, ", %2d", stuckData_memory[38]);
      $fwrite(o, ", %2d", stuckData_memory[39]);
      $fwrite(o, ", %2d", stuckData_memory[40]);
      $fwrite(o, ", %2d", stuckData_memory[41]);
      $fwrite(o, ", %2d", stuckData_memory[42]);
      $fwrite(o, ", %2d", stuckData_memory[43]);
      $fwrite(o, ", %2d", stuckData_memory[44]);
      $fwrite(o, ", %2d", stuckData_memory[45]);
      $fwrite(o, ", %2d", stuckData_memory[46]);
      $fwrite(o, ", %2d", stuckData_memory[47]);
      $fwrite(o, ", %2d", stuckData_memory[48]);
      $fwrite(o, ", %2d", stuckData_memory[49]);
      $fwrite(o, ", %2d", stuckData_memory[50]);
      $fwrite(o, ", %2d", stuckData_memory[51]);
      $fwrite(o, ", %2d", stuckData_memory[52]);
      $fwrite(o, ", %2d", stuckData_memory[53]);
      $fwrite(o, ", %2d", stuckData_memory[54]);
      $fwrite(o, ", %2d", stuckData_memory[55]);
      $fwrite(o, ", %2d", stuckData_memory[56]);
      $fwrite(o, ", %2d", stuckData_memory[57]);
      $fwrite(o, ", %2d", stuckData_memory[58]);
      $fwrite(o, ", %2d", stuckData_memory[59]);
      $fwrite(o, ", %2d", stuckData_memory[60]);
      $fwrite(o, ", %2d", stuckData_memory[61]);
      $fwrite(o, ", %2d", stuckData_memory[62]);
      $fwrite(o, ", %2d", stuckData_memory[63]);
      $fwrite(o, ", %2d", stuckData_memory[64]);
      $fwrite(o, ", %2d", stuckData_memory[65]);
      $fwrite(o, ", %2d", stuckData_memory[66]);
      $fwrite(o, ", %2d", stuckData_memory[67]);
      $fwrite(o, ", %2d", stuckData_memory[68]);
      $fwrite(o, ", %2d", stuckData_memory[69]);
      $fwrite(o, ", %2d", stuckData_memory[70]);
      $fwrite(o, ", %2d", stuckData_memory[71]);
      $fwrite(o, ", %2d", stuckData_memory[72]);
      $fwrite(o, ", %2d", stuckData_memory[73]);
      $fwrite(o, ", %2d", stuckData_memory[74]);
      $fwrite(o, ", %2d", stuckData_memory[75]);
      $fwrite(o, ", %2d", stuckData_memory[76]);
      $fwrite(o, ", %2d", stuckData_memory[77]);
      $fwrite(o, ", %2d", stuckData_memory[78]);
      $fwrite(o, ", %2d", stuckData_memory[79]);
      $fwrite(o, ", %2d", stuckData_memory[80]);
      $fwrite(o, ", %2d", stuckData_memory[81]);
      $fwrite(o, ", %2d", stuckData_memory[82]);
      $fwrite(o, ", %2d", stuckData_memory[83]);
      $fwrite(o, ", %2d", stuckData_memory[84]);
      $fwrite(o, ", %2d", stuckData_memory[85]);
      $fwrite(o, ", %2d", stuckData_memory[86]);
      $fwrite(o, ", %2d", stuckData_memory[87]);
      $fwrite(o, ", %2d", stuckData_memory[88]);
      $fwrite(o, ", %2d", stuckData_memory[89]);
      $fwrite(o, ", %2d", stuckData_memory[90]);
      $fwrite(o, ", %2d", stuckData_memory[91]);
      $fwrite(o, ", %2d", stuckData_memory[92]);
      $fwrite(o, ", %2d", stuckData_memory[93]);
      $fwrite(o, ", %2d", stuckData_memory[94]);
      $fwrite(o, ", %2d", stuckData_memory[95]);
      $fwrite(o, ", %2d", stuckData_memory[96]);
      $fwrite(o, ", %2d", stuckData_memory[97]);
      $fwrite(o, ", %2d", stuckData_memory[98]);
      $fwrite(o, ", %2d", stuckData_memory[99]);
      $fwrite(o, ", %2d", stuckData_memory[100]);
      $fwrite(o, ", %2d", stuckData_memory[101]);
      $fwrite(o, ", %2d", stuckData_memory[102]);
      $fwrite(o, ", %2d", stuckData_memory[103]);
      $fwrite(o, ", %2d", stuckData_memory[104]);
      $fwrite(o, ", %2d", stuckData_memory[105]);
      $fwrite(o, ", %2d", stuckData_memory[106]);
      $fwrite(o, ", %2d", stuckData_memory[107]);
      $fwrite(o, ", %2d", stuckData_memory[108]);
      $fwrite(o, ", %2d", stuckData_memory[109]);
      $fwrite(o, ", %2d", stuckData_memory[110]);
      $fwrite(o, ", %2d", stuckData_memory[111]);
      $fwrite(o, ", %2d", stuckData_memory[112]);
      $fwrite(o, ", %2d", stuckData_memory[113]);
      $fwrite(o, ", %2d", stuckData_memory[114]);
      $fwrite(o, ", %2d", stuckData_memory[115]);
      $fwrite(o, ", %2d", stuckData_memory[116]);
      $fwrite(o, ", %2d", stuckData_memory[117]);
      $fwrite(o, ", %2d", stuckData_memory[118]);
      $fwrite(o, ", %2d", stuckData_memory[119]);
      $fwrite(o, ", %2d", stuckData_memory[120]);
      $fwrite(o, ", %2d", stuckData_memory[121]);
      $fwrite(o, ", %2d", stuckData_memory[122]);
      $fwrite(o, ", %2d", stuckData_memory[123]);
      $fwrite(o, ", %2d", stuckData_memory[124]);
      $fwrite(o, ", %2d", stuckData_memory[125]);
      $fwrite(o, ", %2d", stuckData_memory[126]);
      $fwrite(o, ", %2d", stuckData_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckData_3", stuckData_3_requestedAt, stuckData_3_finishedAt, stuckData_stuckData_3_returnCode, (stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step), (stuckData_3_requestedAt < stuckData_3_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckData_3_index_26", delete_stuckData_3_index_26);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckData_4", stuckData_4_requestedAt, stuckData_4_finishedAt, stuckData_stuckData_4_returnCode, (stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step), (stuckData_4_requestedAt < stuckData_4_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "delete_stuckData_4_index_27", delete_stuckData_4_index_27);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckData_4_value_28", delete_stuckData_4_value_28);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckData_4_value_29", delete_stuckData_4_value_29);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckData_4_value_30", delete_stuckData_4_value_30);

      $fwrite(o, "            %-38s = %1d\n", "delete_stuckData_4_value_31", delete_stuckData_4_value_31);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 6, "delete", 855, delete_pc, delete_returnCode);
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_0", delete_index_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1", delete_size_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_2", delete_isLeaf_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_3", delete_nextFree_3);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_4", delete_Key_0_4);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_5", delete_KeyCompares_0_5);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_6", delete_KeyCollapse_0_6);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_7", delete_Data_0_7);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_8", delete_Key_1_8);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_9", delete_KeyCompares_1_9);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_10", delete_KeyCollapse_1_10);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_11", delete_Data_1_11);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_12", delete_Key_2_12);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_13", delete_KeyCompares_2_13);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_14", delete_KeyCollapse_2_14);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_15", delete_Data_2_15);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_16", delete_Key_3_16);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_17", delete_KeyCompares_3_17);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_18", delete_KeyCollapse_3_18);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_19", delete_Data_3_19);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckKeys_1_index_20", delete_stuckKeys_1_index_20);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckKeys_2_index_21", delete_stuckKeys_2_index_21);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckKeys_2_value_22", delete_stuckKeys_2_value_22);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckKeys_2_value_23", delete_stuckKeys_2_value_23);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckKeys_2_value_24", delete_stuckKeys_2_value_24);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckKeys_2_value_25", delete_stuckKeys_2_value_25);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckData_3_index_26", delete_stuckData_3_index_26);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckData_4_index_27", delete_stuckData_4_index_27);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckData_4_value_28", delete_stuckData_4_value_28);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckData_4_value_29", delete_stuckData_4_value_29);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckData_4_value_30", delete_stuckData_4_value_30);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckData_4_value_31", delete_stuckData_4_value_31);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckSize_5_index_32", delete_stuckSize_5_index_32);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckSize_6_index_33", delete_stuckSize_6_index_33);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckSize_6_value_34", delete_stuckSize_6_value_34);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckIsLeaf_7_index_35", delete_stuckIsLeaf_7_index_35);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckIsLeaf_8_index_36", delete_stuckIsLeaf_8_index_36);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckIsLeaf_8_value_37", delete_stuckIsLeaf_8_value_37);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_38", delete_Found_38);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_39", delete_Key_39);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_40", delete_FoundKey_40);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_41", delete_Data_41);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_42", delete_BtreeIndex_42);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_43", delete_StuckIndex_43);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_44", delete_MergeSuccess_44);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_i_45", delete_i_45);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_k_46", delete_k_46);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_l_47", delete_l_47);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_48", delete_index_48);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_49", delete_size_49);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_50", delete_isLeaf_50);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_51", delete_nextFree_51);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_52", delete_Key_0_52);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_53", delete_KeyCompares_0_53);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_54", delete_KeyCollapse_0_54);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_55", delete_Data_0_55);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_56", delete_Key_1_56);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_57", delete_KeyCompares_1_57);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_58", delete_KeyCollapse_1_58);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_59", delete_Data_1_59);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_60", delete_Key_2_60);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_61", delete_KeyCompares_2_61);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_62", delete_KeyCollapse_2_62);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_63", delete_Data_2_63);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_64", delete_Key_3_64);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_65", delete_KeyCompares_3_65);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_66", delete_KeyCollapse_3_66);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_67", delete_Data_3_67);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_68", delete_Found_68);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_69", delete_Key_69);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_70", delete_FoundKey_70);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_71", delete_Data_71);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_72", delete_BtreeIndex_72);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_73", delete_StuckIndex_73);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_74", delete_MergeSuccess_74);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_75", delete_index_75);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_76", delete_size_76);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_77", delete_isLeaf_77);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_78", delete_nextFree_78);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_79", delete_Key_0_79);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_80", delete_KeyCompares_0_80);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_81", delete_KeyCollapse_0_81);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_82", delete_Data_0_82);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_83", delete_Key_1_83);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_84", delete_KeyCompares_1_84);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_85", delete_KeyCollapse_1_85);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_86", delete_Data_1_86);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_87", delete_Key_2_87);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_88", delete_KeyCompares_2_88);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_89", delete_KeyCollapse_2_89);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_90", delete_Data_2_90);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_91", delete_Key_3_91);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_92", delete_KeyCompares_3_92);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_93", delete_KeyCollapse_3_93);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_94", delete_Data_3_94);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_95", delete_Found_95);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_96", delete_Key_96);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_97", delete_FoundKey_97);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_98", delete_Data_98);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_99", delete_BtreeIndex_99);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_100", delete_StuckIndex_100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_101", delete_MergeSuccess_101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_position_102", delete_position_102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_103", delete_index_103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index1_104", delete_index1_104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_within_105", delete_within_105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_106", delete_isLeaf_106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_107", delete_index_107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_108", delete_size_108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_109", delete_isLeaf_109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_110", delete_nextFree_110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_111", delete_Key_0_111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_112", delete_KeyCompares_0_112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_113", delete_KeyCollapse_0_113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_114", delete_Data_0_114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_115", delete_Key_1_115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_116", delete_KeyCompares_1_116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_117", delete_KeyCollapse_1_117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_118", delete_Data_1_118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_119", delete_Key_2_119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_120", delete_KeyCompares_2_120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_121", delete_KeyCollapse_2_121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_122", delete_Data_2_122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_123", delete_Key_3_123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_124", delete_KeyCompares_3_124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_125", delete_KeyCollapse_3_125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_126", delete_Data_3_126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_127", delete_Found_127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_128", delete_Key_128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_129", delete_FoundKey_129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_130", delete_Data_130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_131", delete_BtreeIndex_131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_132", delete_StuckIndex_132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_133", delete_MergeSuccess_133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_134", delete_index_134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_135", delete_size_135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_136", delete_isLeaf_136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_137", delete_nextFree_137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_138", delete_Key_0_138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_139", delete_KeyCompares_0_139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_140", delete_KeyCollapse_0_140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_141", delete_Data_0_141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_142", delete_Key_1_142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_143", delete_KeyCompares_1_143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_144", delete_KeyCollapse_1_144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_145", delete_Data_1_145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_146", delete_Key_2_146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_147", delete_KeyCompares_2_147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_148", delete_KeyCollapse_2_148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_149", delete_Data_2_149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_150", delete_Key_3_150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_151", delete_KeyCompares_3_151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_152", delete_KeyCollapse_3_152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_153", delete_Data_3_153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_154", delete_Found_154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_155", delete_Key_155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_156", delete_FoundKey_156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_157", delete_Data_157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_158", delete_BtreeIndex_158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_159", delete_StuckIndex_159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_160", delete_MergeSuccess_160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_161", delete_index_161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_162", delete_size_162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_163", delete_isLeaf_163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_164", delete_nextFree_164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_165", delete_Key_0_165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_166", delete_KeyCompares_0_166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_167", delete_KeyCollapse_0_167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_168", delete_Data_0_168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_169", delete_Key_1_169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_170", delete_KeyCompares_1_170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_171", delete_KeyCollapse_1_171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_172", delete_Data_1_172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_173", delete_Key_2_173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_174", delete_KeyCompares_2_174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_175", delete_KeyCollapse_2_175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_176", delete_Data_2_176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_177", delete_Key_3_177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_178", delete_KeyCompares_3_178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_179", delete_KeyCollapse_3_179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_180", delete_Data_3_180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_181", delete_Found_181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_182", delete_Key_182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_183", delete_FoundKey_183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_184", delete_Data_184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_185", delete_BtreeIndex_185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_186", delete_StuckIndex_186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_187", delete_MergeSuccess_187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_188", delete_childKey_188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_189", delete_childData_189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_190", delete_indexLeft_190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_191", delete_indexRight_191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_192", delete_midKey_192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_193", delete_success_193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_194", delete_test_194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_195", delete_next_195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_freeNext_9_index_196", delete_freeNext_9_index_196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_freeNext_10_index_197", delete_freeNext_10_index_197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_freeNext_10_value_198", delete_freeNext_10_value_198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckIsFree_11_index_199", delete_stuckIsFree_11_index_199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_stuckIsFree_11_value_200", delete_stuckIsFree_11_value_200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_201", delete_root_201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_202", delete_isFree_202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_203", delete_next_203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_204", delete_root_204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_205", delete_isFree_205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_206", delete_index_206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_207", delete_size_207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_208", delete_isLeaf_208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_209", delete_nextFree_209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_210", delete_Key_0_210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_211", delete_KeyCompares_0_211);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_212", delete_KeyCollapse_0_212);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_213", delete_Data_0_213);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_214", delete_Key_1_214);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_215", delete_KeyCompares_1_215);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_216", delete_KeyCollapse_1_216);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_217", delete_Data_1_217);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_218", delete_Key_2_218);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_219", delete_KeyCompares_2_219);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_220", delete_KeyCollapse_2_220);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_221", delete_Data_2_221);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_222", delete_Key_3_222);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_223", delete_KeyCompares_3_223);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_224", delete_KeyCollapse_3_224);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_225", delete_Data_3_225);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_226", delete_Found_226);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_227", delete_Key_227);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_228", delete_FoundKey_228);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_229", delete_Data_229);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_230", delete_BtreeIndex_230);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_231", delete_StuckIndex_231);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_232", delete_MergeSuccess_232);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_233", delete_index_233);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_234", delete_size_234);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_235", delete_isLeaf_235);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_236", delete_nextFree_236);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_237", delete_Key_0_237);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_238", delete_KeyCompares_0_238);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_239", delete_KeyCollapse_0_239);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_240", delete_Data_0_240);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_241", delete_Key_1_241);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_242", delete_KeyCompares_1_242);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_243", delete_KeyCollapse_1_243);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_244", delete_Data_1_244);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_245", delete_Key_2_245);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_246", delete_KeyCompares_2_246);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_247", delete_KeyCollapse_2_247);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_248", delete_Data_2_248);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_249", delete_Key_3_249);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_250", delete_KeyCompares_3_250);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_251", delete_KeyCollapse_3_251);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_252", delete_Data_3_252);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_253", delete_Found_253);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_254", delete_Key_254);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_255", delete_FoundKey_255);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_256", delete_Data_256);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_257", delete_BtreeIndex_257);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_258", delete_StuckIndex_258);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_259", delete_MergeSuccess_259);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_260", delete_index_260);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_261", delete_size_261);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_262", delete_isLeaf_262);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_263", delete_nextFree_263);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_264", delete_Key_0_264);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_265", delete_KeyCompares_0_265);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_266", delete_KeyCollapse_0_266);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_267", delete_Data_0_267);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_268", delete_Key_1_268);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_269", delete_KeyCompares_1_269);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_270", delete_KeyCollapse_1_270);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_271", delete_Data_1_271);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_272", delete_Key_2_272);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_273", delete_KeyCompares_2_273);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_274", delete_KeyCollapse_2_274);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_275", delete_Data_2_275);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_276", delete_Key_3_276);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_277", delete_KeyCompares_3_277);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_278", delete_KeyCollapse_3_278);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_279", delete_Data_3_279);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_280", delete_Found_280);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_281", delete_Key_281);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_282", delete_FoundKey_282);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_283", delete_Data_283);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_284", delete_BtreeIndex_284);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_285", delete_StuckIndex_285);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_286", delete_MergeSuccess_286);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_287", delete_childKey_287);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_288", delete_leftChild_288);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_289", delete_rightChild_289);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_290", delete_childData_290);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_291", delete_indexLeft_291);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_292", delete_indexRight_292);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_293", delete_midKey_293);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_294", delete_success_294);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_295", delete_test_295);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_296", delete_next_296);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_297", delete_root_297);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_298", delete_isFree_298);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_299", delete_next_299);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_300", delete_root_300);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_301", delete_isFree_301);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_302", delete_index_302);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_303", delete_size_303);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_304", delete_isLeaf_304);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_305", delete_nextFree_305);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_306", delete_Key_0_306);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_307", delete_KeyCompares_0_307);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_308", delete_KeyCollapse_0_308);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_309", delete_Data_0_309);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_310", delete_Key_1_310);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_311", delete_KeyCompares_1_311);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_312", delete_KeyCollapse_1_312);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_313", delete_Data_1_313);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_314", delete_Key_2_314);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_315", delete_KeyCompares_2_315);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_316", delete_KeyCollapse_2_316);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_317", delete_Data_2_317);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_318", delete_Key_3_318);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_319", delete_KeyCompares_3_319);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_320", delete_KeyCollapse_3_320);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_321", delete_Data_3_321);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_322", delete_Found_322);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_323", delete_Key_323);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_324", delete_FoundKey_324);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_325", delete_Data_325);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_326", delete_BtreeIndex_326);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_327", delete_StuckIndex_327);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_328", delete_MergeSuccess_328);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_329", delete_index_329);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_330", delete_size_330);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_331", delete_isLeaf_331);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_332", delete_nextFree_332);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_333", delete_Key_0_333);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_334", delete_KeyCompares_0_334);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_335", delete_KeyCollapse_0_335);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_336", delete_Data_0_336);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_337", delete_Key_1_337);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_338", delete_KeyCompares_1_338);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_339", delete_KeyCollapse_1_339);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_340", delete_Data_1_340);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_341", delete_Key_2_341);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_342", delete_KeyCompares_2_342);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_343", delete_KeyCollapse_2_343);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_344", delete_Data_2_344);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_345", delete_Key_3_345);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_346", delete_KeyCompares_3_346);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_347", delete_KeyCollapse_3_347);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_348", delete_Data_3_348);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_349", delete_Found_349);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_350", delete_Key_350);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_351", delete_FoundKey_351);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_352", delete_Data_352);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_353", delete_BtreeIndex_353);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_354", delete_StuckIndex_354);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_355", delete_MergeSuccess_355);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_356", delete_childKey_356);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_357", delete_size_357);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_358", delete_childData_358);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_359", delete_indexLeft_359);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_360", delete_indexRight_360);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_361", delete_midKey_361);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_362", delete_success_362);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_363", delete_test_363);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_364", delete_next_364);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_365", delete_root_365);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_366", delete_isFree_366);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_367", delete_index_367);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_368", delete_size_368);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_369", delete_isLeaf_369);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_370", delete_nextFree_370);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_371", delete_Key_0_371);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_372", delete_KeyCompares_0_372);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_373", delete_KeyCollapse_0_373);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_374", delete_Data_0_374);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_375", delete_Key_1_375);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_376", delete_KeyCompares_1_376);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_377", delete_KeyCollapse_1_377);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_378", delete_Data_1_378);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_379", delete_Key_2_379);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_380", delete_KeyCompares_2_380);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_381", delete_KeyCollapse_2_381);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_382", delete_Data_2_382);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_383", delete_Key_3_383);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_384", delete_KeyCompares_3_384);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_385", delete_KeyCollapse_3_385);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_386", delete_Data_3_386);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_387", delete_Found_387);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_388", delete_Key_388);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_389", delete_FoundKey_389);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_390", delete_Data_390);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_391", delete_BtreeIndex_391);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_392", delete_StuckIndex_392);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_393", delete_MergeSuccess_393);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_394", delete_index_394);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_395", delete_size_395);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_396", delete_isLeaf_396);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_397", delete_nextFree_397);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_398", delete_Key_0_398);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_399", delete_KeyCompares_0_399);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_400", delete_KeyCollapse_0_400);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_401", delete_Data_0_401);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_402", delete_Key_1_402);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_403", delete_KeyCompares_1_403);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_404", delete_KeyCollapse_1_404);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_405", delete_Data_1_405);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_406", delete_Key_2_406);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_407", delete_KeyCompares_2_407);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_408", delete_KeyCollapse_2_408);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_409", delete_Data_2_409);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_410", delete_Key_3_410);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_411", delete_KeyCompares_3_411);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_412", delete_KeyCollapse_3_412);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_413", delete_Data_3_413);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_414", delete_Found_414);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_415", delete_Key_415);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_416", delete_FoundKey_416);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_417", delete_Data_417);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_418", delete_BtreeIndex_418);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_419", delete_StuckIndex_419);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_420", delete_MergeSuccess_420);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_421", delete_childKey_421);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_422", delete_size_422);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_423", delete_childData_423);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_424", delete_indexLeft_424);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_425", delete_indexRight_425);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_426", delete_midKey_426);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_427", delete_success_427);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_428", delete_test_428);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_429", delete_next_429);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_430", delete_root_430);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_431", delete_isFree_431);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_432", delete_index_432);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_433", delete_size_433);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_434", delete_isLeaf_434);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_435", delete_nextFree_435);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_436", delete_Key_0_436);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_437", delete_KeyCompares_0_437);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_438", delete_KeyCollapse_0_438);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_439", delete_Data_0_439);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_440", delete_Key_1_440);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_441", delete_KeyCompares_1_441);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_442", delete_KeyCollapse_1_442);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_443", delete_Data_1_443);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_444", delete_Key_2_444);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_445", delete_KeyCompares_2_445);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_446", delete_KeyCollapse_2_446);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_447", delete_Data_2_447);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_448", delete_Key_3_448);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_449", delete_KeyCompares_3_449);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_450", delete_KeyCollapse_3_450);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_451", delete_Data_3_451);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_452", delete_Found_452);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_453", delete_Key_453);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_454", delete_FoundKey_454);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_455", delete_Data_455);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_456", delete_BtreeIndex_456);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_457", delete_StuckIndex_457);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_458", delete_MergeSuccess_458);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_459", delete_index_459);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_460", delete_size_460);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_461", delete_isLeaf_461);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_462", delete_nextFree_462);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_463", delete_Key_0_463);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_464", delete_KeyCompares_0_464);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_465", delete_KeyCollapse_0_465);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_466", delete_Data_0_466);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_467", delete_Key_1_467);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_468", delete_KeyCompares_1_468);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_469", delete_KeyCollapse_1_469);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_470", delete_Data_1_470);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_471", delete_Key_2_471);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_472", delete_KeyCompares_2_472);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_473", delete_KeyCollapse_2_473);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_474", delete_Data_2_474);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_475", delete_Key_3_475);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_476", delete_KeyCompares_3_476);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_477", delete_KeyCollapse_3_477);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_478", delete_Data_3_478);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_479", delete_Found_479);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_480", delete_Key_480);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_481", delete_FoundKey_481);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_482", delete_Data_482);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_483", delete_BtreeIndex_483);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_484", delete_StuckIndex_484);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_485", delete_MergeSuccess_485);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_486", delete_childKey_486);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_487", delete_childData_487);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_488", delete_indexLeft_488);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_489", delete_indexRight_489);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_490", delete_midKey_490);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_491", delete_success_491);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_492", delete_test_492);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_493", delete_next_493);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_494", delete_root_494);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_495", delete_isFree_495);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_496", delete_index_496);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_497", delete_size_497);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_498", delete_isLeaf_498);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_499", delete_nextFree_499);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_500", delete_Key_0_500);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_501", delete_KeyCompares_0_501);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_502", delete_KeyCollapse_0_502);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_503", delete_Data_0_503);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_504", delete_Key_1_504);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_505", delete_KeyCompares_1_505);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_506", delete_KeyCollapse_1_506);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_507", delete_Data_1_507);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_508", delete_Key_2_508);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_509", delete_KeyCompares_2_509);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_510", delete_KeyCollapse_2_510);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_511", delete_Data_2_511);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_512", delete_Key_3_512);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_513", delete_KeyCompares_3_513);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_514", delete_KeyCollapse_3_514);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_515", delete_Data_3_515);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_516", delete_Found_516);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_517", delete_Key_517);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_518", delete_FoundKey_518);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_519", delete_Data_519);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_520", delete_BtreeIndex_520);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_521", delete_StuckIndex_521);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_522", delete_MergeSuccess_522);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_523", delete_index_523);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_524", delete_size_524);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_525", delete_isLeaf_525);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_526", delete_nextFree_526);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_527", delete_Key_0_527);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_528", delete_KeyCompares_0_528);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_529", delete_KeyCollapse_0_529);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_530", delete_Data_0_530);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_531", delete_Key_1_531);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_532", delete_KeyCompares_1_532);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_533", delete_KeyCollapse_1_533);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_534", delete_Data_1_534);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_535", delete_Key_2_535);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_536", delete_KeyCompares_2_536);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_537", delete_KeyCollapse_2_537);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_538", delete_Data_2_538);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_539", delete_Key_3_539);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_540", delete_KeyCompares_3_540);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_541", delete_KeyCollapse_3_541);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_542", delete_Data_3_542);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_543", delete_Found_543);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_544", delete_Key_544);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_545", delete_FoundKey_545);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_546", delete_Data_546);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_547", delete_BtreeIndex_547);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_548", delete_StuckIndex_548);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_549", delete_MergeSuccess_549);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_550", delete_childKey_550);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_551", delete_leftChild_551);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_552", delete_rightChild_552);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_553", delete_childData_553);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_554", delete_indexLeft_554);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_555", delete_indexRight_555);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_556", delete_midKey_556);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_557", delete_success_557);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_558", delete_test_558);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_559", delete_next_559);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_560", delete_root_560);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_561", delete_isFree_561);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_562", delete_index_562);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_563", delete_size_563);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_564", delete_isLeaf_564);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_565", delete_nextFree_565);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_566", delete_Key_0_566);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_567", delete_KeyCompares_0_567);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_568", delete_KeyCollapse_0_568);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_569", delete_Data_0_569);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_570", delete_Key_1_570);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_571", delete_KeyCompares_1_571);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_572", delete_KeyCollapse_1_572);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_573", delete_Data_1_573);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_574", delete_Key_2_574);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_575", delete_KeyCompares_2_575);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_576", delete_KeyCollapse_2_576);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_577", delete_Data_2_577);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_578", delete_Key_3_578);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_579", delete_KeyCompares_3_579);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_580", delete_KeyCollapse_3_580);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_581", delete_Data_3_581);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_582", delete_Found_582);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_583", delete_Key_583);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_584", delete_FoundKey_584);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_585", delete_Data_585);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_586", delete_BtreeIndex_586);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_587", delete_StuckIndex_587);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_588", delete_MergeSuccess_588);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_589", delete_index_589);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_590", delete_size_590);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_591", delete_isLeaf_591);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_592", delete_nextFree_592);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_593", delete_Key_0_593);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_594", delete_KeyCompares_0_594);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_595", delete_KeyCollapse_0_595);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_596", delete_Data_0_596);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_597", delete_Key_1_597);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_598", delete_KeyCompares_1_598);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_599", delete_KeyCollapse_1_599);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_600", delete_Data_1_600);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_601", delete_Key_2_601);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_602", delete_KeyCompares_2_602);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_603", delete_KeyCollapse_2_603);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_604", delete_Data_2_604);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_605", delete_Key_3_605);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_606", delete_KeyCompares_3_606);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_607", delete_KeyCollapse_3_607);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_608", delete_Data_3_608);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_609", delete_Found_609);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_610", delete_Key_610);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_611", delete_FoundKey_611);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_612", delete_Data_612);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_613", delete_BtreeIndex_613);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_614", delete_StuckIndex_614);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_615", delete_MergeSuccess_615);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_616", delete_childKey_616);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_617", delete_childData_617);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_618", delete_indexLeft_618);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_619", delete_indexRight_619);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_620", delete_midKey_620);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_621", delete_success_621);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_622", delete_test_622);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_623", delete_next_623);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_624", delete_root_624);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_625", delete_isFree_625);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_626", delete_index_626);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_627", delete_size_627);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_628", delete_isLeaf_628);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_629", delete_nextFree_629);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_630", delete_Key_0_630);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_631", delete_KeyCompares_0_631);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_632", delete_KeyCollapse_0_632);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_633", delete_Data_0_633);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_634", delete_Key_1_634);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_635", delete_KeyCompares_1_635);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_636", delete_KeyCollapse_1_636);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_637", delete_Data_1_637);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_638", delete_Key_2_638);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_639", delete_KeyCompares_2_639);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_640", delete_KeyCollapse_2_640);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_641", delete_Data_2_641);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_642", delete_Key_3_642);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_643", delete_KeyCompares_3_643);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_644", delete_KeyCollapse_3_644);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_645", delete_Data_3_645);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_646", delete_Found_646);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_647", delete_Key_647);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_648", delete_FoundKey_648);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_649", delete_Data_649);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_650", delete_BtreeIndex_650);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_651", delete_StuckIndex_651);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_652", delete_MergeSuccess_652);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_653", delete_index_653);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_654", delete_size_654);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_655", delete_isLeaf_655);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_656", delete_nextFree_656);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_657", delete_Key_0_657);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_658", delete_KeyCompares_0_658);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_659", delete_KeyCollapse_0_659);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_660", delete_Data_0_660);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_661", delete_Key_1_661);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_662", delete_KeyCompares_1_662);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_663", delete_KeyCollapse_1_663);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_664", delete_Data_1_664);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_665", delete_Key_2_665);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_666", delete_KeyCompares_2_666);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_667", delete_KeyCollapse_2_667);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_668", delete_Data_2_668);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_669", delete_Key_3_669);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_670", delete_KeyCompares_3_670);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_671", delete_KeyCollapse_3_671);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_672", delete_Data_3_672);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_673", delete_Found_673);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_674", delete_Key_674);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_675", delete_FoundKey_675);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_676", delete_Data_676);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_677", delete_BtreeIndex_677);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_678", delete_StuckIndex_678);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_679", delete_MergeSuccess_679);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_680", delete_childKey_680);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_681", delete_leftChild_681);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_682", delete_rightChild_682);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_683", delete_childData_683);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_684", delete_indexLeft_684);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_685", delete_indexRight_685);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_686", delete_midKey_686);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_687", delete_success_687);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_688", delete_test_688);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_689", delete_next_689);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_690", delete_root_690);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_691", delete_isFree_691);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_692", delete_index_692);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_693", delete_size_693);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_694", delete_isLeaf_694);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_695", delete_nextFree_695);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_696", delete_Key_0_696);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_697", delete_KeyCompares_0_697);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_698", delete_KeyCollapse_0_698);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_699", delete_Data_0_699);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_700", delete_Key_1_700);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_701", delete_KeyCompares_1_701);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_702", delete_KeyCollapse_1_702);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_703", delete_Data_1_703);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_704", delete_Key_2_704);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_705", delete_KeyCompares_2_705);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_706", delete_KeyCollapse_2_706);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_707", delete_Data_2_707);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_708", delete_Key_3_708);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_709", delete_KeyCompares_3_709);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_710", delete_KeyCollapse_3_710);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_711", delete_Data_3_711);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_712", delete_Found_712);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_713", delete_Key_713);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_714", delete_FoundKey_714);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_715", delete_Data_715);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_716", delete_BtreeIndex_716);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_717", delete_StuckIndex_717);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_718", delete_MergeSuccess_718);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_719", delete_index_719);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_720", delete_size_720);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_721", delete_isLeaf_721);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_722", delete_nextFree_722);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_723", delete_Key_0_723);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_724", delete_KeyCompares_0_724);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_725", delete_KeyCollapse_0_725);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_726", delete_Data_0_726);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_727", delete_Key_1_727);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_728", delete_KeyCompares_1_728);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_729", delete_KeyCollapse_1_729);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_730", delete_Data_1_730);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_731", delete_Key_2_731);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_732", delete_KeyCompares_2_732);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_733", delete_KeyCollapse_2_733);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_734", delete_Data_2_734);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_735", delete_Key_3_735);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_736", delete_KeyCompares_3_736);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_737", delete_KeyCollapse_3_737);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_738", delete_Data_3_738);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_739", delete_Found_739);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_740", delete_Key_740);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_741", delete_FoundKey_741);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_742", delete_Data_742);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_743", delete_BtreeIndex_743);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_744", delete_StuckIndex_744);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_745", delete_MergeSuccess_745);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_746", delete_childKey_746);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_747", delete_childData_747);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_748", delete_indexLeft_748);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_749", delete_indexRight_749);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_750", delete_midKey_750);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_751", delete_success_751);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_752", delete_test_752);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_753", delete_next_753);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_754", delete_root_754);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_755", delete_isFree_755);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_756", delete_index_756);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_757", delete_size_757);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_758", delete_isLeaf_758);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_759", delete_nextFree_759);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_760", delete_Key_0_760);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_761", delete_KeyCompares_0_761);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_762", delete_KeyCollapse_0_762);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_763", delete_Data_0_763);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_764", delete_Key_1_764);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_765", delete_KeyCompares_1_765);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_766", delete_KeyCollapse_1_766);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_767", delete_Data_1_767);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_768", delete_Key_2_768);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_769", delete_KeyCompares_2_769);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_770", delete_KeyCollapse_2_770);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_771", delete_Data_2_771);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_772", delete_Key_3_772);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_773", delete_KeyCompares_3_773);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_774", delete_KeyCollapse_3_774);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_775", delete_Data_3_775);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_776", delete_Found_776);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_777", delete_Key_777);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_778", delete_FoundKey_778);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_779", delete_Data_779);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_780", delete_BtreeIndex_780);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_781", delete_StuckIndex_781);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_782", delete_MergeSuccess_782);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_783", delete_index_783);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_784", delete_size_784);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_785", delete_isLeaf_785);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_786", delete_nextFree_786);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_787", delete_Key_0_787);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_788", delete_KeyCompares_0_788);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_789", delete_KeyCollapse_0_789);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_790", delete_Data_0_790);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_791", delete_Key_1_791);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_792", delete_KeyCompares_1_792);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_793", delete_KeyCollapse_1_793);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_794", delete_Data_1_794);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_795", delete_Key_2_795);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_796", delete_KeyCompares_2_796);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_797", delete_KeyCollapse_2_797);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_798", delete_Data_2_798);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_799", delete_Key_3_799);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_800", delete_KeyCompares_3_800);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_801", delete_KeyCollapse_3_801);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_802", delete_Data_3_802);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_803", delete_Found_803);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_804", delete_Key_804);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_805", delete_FoundKey_805);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_806", delete_Data_806);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_807", delete_BtreeIndex_807);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_808", delete_StuckIndex_808);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_809", delete_MergeSuccess_809);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_810", delete_childKey_810);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_811", delete_leftChild_811);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_812", delete_rightChild_812);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_813", delete_childData_813);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_814", delete_indexLeft_814);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_815", delete_indexRight_815);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_816", delete_midKey_816);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_817", delete_success_817);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_818", delete_test_818);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_819", delete_next_819);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_820", delete_root_820);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_821", delete_isFree_821);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_822", delete_index_822);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_823", delete_size_823);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_824", delete_isLeaf_824);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_825", delete_nextFree_825);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_826", delete_Key_0_826);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_827", delete_KeyCompares_0_827);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_828", delete_KeyCollapse_0_828);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_829", delete_Data_0_829);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_830", delete_Key_1_830);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_831", delete_KeyCompares_1_831);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_832", delete_KeyCollapse_1_832);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_833", delete_Data_1_833);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_834", delete_Key_2_834);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_835", delete_KeyCompares_2_835);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_836", delete_KeyCollapse_2_836);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_837", delete_Data_2_837);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_838", delete_Key_3_838);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_839", delete_KeyCompares_3_839);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_840", delete_KeyCollapse_3_840);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_841", delete_Data_3_841);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_842", delete_Found_842);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_843", delete_Key_843);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_844", delete_FoundKey_844);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_845", delete_Data_845);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_846", delete_BtreeIndex_846);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_847", delete_StuckIndex_847);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_848", delete_MergeSuccess_848);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_849", delete_index_849);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_850", delete_size_850);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_851", delete_isLeaf_851);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_852", delete_nextFree_852);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_853", delete_Key_0_853);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_854", delete_KeyCompares_0_854);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_855", delete_KeyCollapse_0_855);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_856", delete_Data_0_856);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_857", delete_Key_1_857);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_858", delete_KeyCompares_1_858);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_859", delete_KeyCollapse_1_859);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_860", delete_Data_1_860);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_861", delete_Key_2_861);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_862", delete_KeyCompares_2_862);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_863", delete_KeyCollapse_2_863);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_864", delete_Data_2_864);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_865", delete_Key_3_865);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_866", delete_KeyCompares_3_866);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_867", delete_KeyCollapse_3_867);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_868", delete_Data_3_868);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_869", delete_Found_869);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_870", delete_Key_870);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_871", delete_FoundKey_871);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_872", delete_Data_872);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_873", delete_BtreeIndex_873);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_874", delete_StuckIndex_874);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_875", delete_MergeSuccess_875);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_876", delete_childKey_876);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_877", delete_childData_877);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_878", delete_indexLeft_878);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_879", delete_indexRight_879);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_880", delete_midKey_880);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_881", delete_success_881);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_882", delete_test_882);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_883", delete_next_883);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_884", delete_root_884);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_885", delete_isFree_885);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_886", delete_index_886);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_887", delete_size_887);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_888", delete_isLeaf_888);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_889", delete_nextFree_889);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_890", delete_Key_0_890);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_891", delete_KeyCompares_0_891);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_892", delete_KeyCollapse_0_892);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_893", delete_Data_0_893);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_894", delete_Key_1_894);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_895", delete_KeyCompares_1_895);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_896", delete_KeyCollapse_1_896);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_897", delete_Data_1_897);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_898", delete_Key_2_898);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_899", delete_KeyCompares_2_899);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_900", delete_KeyCollapse_2_900);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_901", delete_Data_2_901);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_902", delete_Key_3_902);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_903", delete_KeyCompares_3_903);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_904", delete_KeyCollapse_3_904);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_905", delete_Data_3_905);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_906", delete_Found_906);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_907", delete_Key_907);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_908", delete_FoundKey_908);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_909", delete_Data_909);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_910", delete_BtreeIndex_910);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_911", delete_StuckIndex_911);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_912", delete_MergeSuccess_912);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_913", delete_index_913);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_914", delete_size_914);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_915", delete_isLeaf_915);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_916", delete_nextFree_916);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_917", delete_Key_0_917);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_918", delete_KeyCompares_0_918);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_919", delete_KeyCollapse_0_919);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_920", delete_Data_0_920);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_921", delete_Key_1_921);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_922", delete_KeyCompares_1_922);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_923", delete_KeyCollapse_1_923);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_924", delete_Data_1_924);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_925", delete_Key_2_925);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_926", delete_KeyCompares_2_926);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_927", delete_KeyCollapse_2_927);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_928", delete_Data_2_928);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_929", delete_Key_3_929);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_930", delete_KeyCompares_3_930);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_931", delete_KeyCollapse_3_931);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_932", delete_Data_3_932);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_933", delete_Found_933);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_934", delete_Key_934);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_935", delete_FoundKey_935);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_936", delete_Data_936);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_937", delete_BtreeIndex_937);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_938", delete_StuckIndex_938);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_939", delete_MergeSuccess_939);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_940", delete_childKey_940);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_941", delete_leftChild_941);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_942", delete_rightChild_942);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_943", delete_childData_943);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_944", delete_indexLeft_944);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_945", delete_indexRight_945);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_946", delete_midKey_946);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_947", delete_success_947);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_948", delete_test_948);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_949", delete_next_949);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_950", delete_root_950);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_951", delete_isFree_951);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_952", delete_index_952);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_953", delete_size_953);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_954", delete_isLeaf_954);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_955", delete_nextFree_955);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_956", delete_Key_0_956);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_957", delete_KeyCompares_0_957);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_958", delete_KeyCollapse_0_958);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_959", delete_Data_0_959);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_960", delete_Key_1_960);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_961", delete_KeyCompares_1_961);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_962", delete_KeyCollapse_1_962);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_963", delete_Data_1_963);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_964", delete_Key_2_964);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_965", delete_KeyCompares_2_965);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_966", delete_KeyCollapse_2_966);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_967", delete_Data_2_967);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_968", delete_Key_3_968);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_969", delete_KeyCompares_3_969);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_970", delete_KeyCollapse_3_970);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_971", delete_Data_3_971);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_972", delete_Found_972);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_973", delete_Key_973);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_974", delete_FoundKey_974);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_975", delete_Data_975);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_976", delete_BtreeIndex_976);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_977", delete_StuckIndex_977);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_978", delete_MergeSuccess_978);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_979", delete_index_979);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_980", delete_size_980);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_981", delete_isLeaf_981);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_982", delete_nextFree_982);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_983", delete_Key_0_983);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_984", delete_KeyCompares_0_984);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_985", delete_KeyCollapse_0_985);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_986", delete_Data_0_986);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_987", delete_Key_1_987);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_988", delete_KeyCompares_1_988);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_989", delete_KeyCollapse_1_989);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_990", delete_Data_1_990);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_991", delete_Key_2_991);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_992", delete_KeyCompares_2_992);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_993", delete_KeyCollapse_2_993);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_994", delete_Data_2_994);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_995", delete_Key_3_995);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_996", delete_KeyCompares_3_996);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_997", delete_KeyCollapse_3_997);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_998", delete_Data_3_998);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_999", delete_Found_999);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1000", delete_Key_1000);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1001", delete_FoundKey_1001);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1002", delete_Data_1002);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1003", delete_BtreeIndex_1003);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1004", delete_StuckIndex_1004);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1005", delete_MergeSuccess_1005);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_1006", delete_childKey_1006);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_1007", delete_childData_1007);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_1008", delete_indexLeft_1008);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_1009", delete_indexRight_1009);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_1010", delete_midKey_1010);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_1011", delete_success_1011);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_1012", delete_test_1012);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_1013", delete_next_1013);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_1014", delete_root_1014);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_1015", delete_isFree_1015);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_1016", delete_index_1016);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1017", delete_size_1017);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_1018", delete_isLeaf_1018);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_1019", delete_nextFree_1019);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_1020", delete_Key_0_1020);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_1021", delete_KeyCompares_0_1021);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_1022", delete_KeyCollapse_0_1022);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_1023", delete_Data_0_1023);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_1024", delete_Key_1_1024);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_1025", delete_KeyCompares_1_1025);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_1026", delete_KeyCollapse_1_1026);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_1027", delete_Data_1_1027);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_1028", delete_Key_2_1028);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_1029", delete_KeyCompares_2_1029);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_1030", delete_KeyCollapse_2_1030);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_1031", delete_Data_2_1031);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_1032", delete_Key_3_1032);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_1033", delete_KeyCompares_3_1033);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_1034", delete_KeyCollapse_3_1034);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_1035", delete_Data_3_1035);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_1036", delete_Found_1036);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1037", delete_Key_1037);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1038", delete_FoundKey_1038);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1039", delete_Data_1039);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1040", delete_BtreeIndex_1040);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1041", delete_StuckIndex_1041);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1042", delete_MergeSuccess_1042);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_1043", delete_index_1043);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1044", delete_size_1044);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_1045", delete_isLeaf_1045);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_1046", delete_nextFree_1046);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_1047", delete_Key_0_1047);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_1048", delete_KeyCompares_0_1048);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_1049", delete_KeyCollapse_0_1049);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_1050", delete_Data_0_1050);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_1051", delete_Key_1_1051);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_1052", delete_KeyCompares_1_1052);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_1053", delete_KeyCollapse_1_1053);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_1054", delete_Data_1_1054);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_1055", delete_Key_2_1055);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_1056", delete_KeyCompares_2_1056);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_1057", delete_KeyCollapse_2_1057);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_1058", delete_Data_2_1058);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_1059", delete_Key_3_1059);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_1060", delete_KeyCompares_3_1060);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_1061", delete_KeyCollapse_3_1061);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_1062", delete_Data_3_1062);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_1063", delete_Found_1063);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1064", delete_Key_1064);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1065", delete_FoundKey_1065);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1066", delete_Data_1066);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1067", delete_BtreeIndex_1067);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1068", delete_StuckIndex_1068);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1069", delete_MergeSuccess_1069);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_1070", delete_childKey_1070);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_1071", delete_leftChild_1071);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_1072", delete_rightChild_1072);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_1073", delete_childData_1073);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_1074", delete_indexLeft_1074);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_1075", delete_indexRight_1075);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_1076", delete_midKey_1076);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_1077", delete_success_1077);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_1078", delete_test_1078);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_1079", delete_next_1079);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_1080", delete_root_1080);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_1081", delete_isFree_1081);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_1082", delete_index_1082);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1083", delete_size_1083);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_1084", delete_isLeaf_1084);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_1085", delete_nextFree_1085);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_1086", delete_Key_0_1086);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_1087", delete_KeyCompares_0_1087);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_1088", delete_KeyCollapse_0_1088);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_1089", delete_Data_0_1089);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_1090", delete_Key_1_1090);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_1091", delete_KeyCompares_1_1091);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_1092", delete_KeyCollapse_1_1092);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_1093", delete_Data_1_1093);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_1094", delete_Key_2_1094);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_1095", delete_KeyCompares_2_1095);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_1096", delete_KeyCollapse_2_1096);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_1097", delete_Data_2_1097);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_1098", delete_Key_3_1098);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_1099", delete_KeyCompares_3_1099);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_1100", delete_KeyCollapse_3_1100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_1101", delete_Data_3_1101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_1102", delete_Found_1102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1103", delete_Key_1103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1104", delete_FoundKey_1104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1105", delete_Data_1105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1106", delete_BtreeIndex_1106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1107", delete_StuckIndex_1107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1108", delete_MergeSuccess_1108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_1109", delete_index_1109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1110", delete_size_1110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_1111", delete_isLeaf_1111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_1112", delete_nextFree_1112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_1113", delete_Key_0_1113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_1114", delete_KeyCompares_0_1114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_1115", delete_KeyCollapse_0_1115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_1116", delete_Data_0_1116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_1117", delete_Key_1_1117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_1118", delete_KeyCompares_1_1118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_1119", delete_KeyCollapse_1_1119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_1120", delete_Data_1_1120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_1121", delete_Key_2_1121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_1122", delete_KeyCompares_2_1122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_1123", delete_KeyCollapse_2_1123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_1124", delete_Data_2_1124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_1125", delete_Key_3_1125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_1126", delete_KeyCompares_3_1126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_1127", delete_KeyCollapse_3_1127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_1128", delete_Data_3_1128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_1129", delete_Found_1129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1130", delete_Key_1130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1131", delete_FoundKey_1131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1132", delete_Data_1132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1133", delete_BtreeIndex_1133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1134", delete_StuckIndex_1134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1135", delete_MergeSuccess_1135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_1136", delete_childKey_1136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_1137", delete_childData_1137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_1138", delete_indexLeft_1138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_1139", delete_indexRight_1139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_1140", delete_midKey_1140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_1141", delete_success_1141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_1142", delete_test_1142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_1143", delete_next_1143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_1144", delete_root_1144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_1145", delete_isFree_1145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_1146", delete_index_1146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1147", delete_size_1147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_1148", delete_isLeaf_1148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_1149", delete_nextFree_1149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_1150", delete_Key_0_1150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_1151", delete_KeyCompares_0_1151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_1152", delete_KeyCollapse_0_1152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_1153", delete_Data_0_1153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_1154", delete_Key_1_1154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_1155", delete_KeyCompares_1_1155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_1156", delete_KeyCollapse_1_1156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_1157", delete_Data_1_1157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_1158", delete_Key_2_1158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_1159", delete_KeyCompares_2_1159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_1160", delete_KeyCollapse_2_1160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_1161", delete_Data_2_1161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_1162", delete_Key_3_1162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_1163", delete_KeyCompares_3_1163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_1164", delete_KeyCollapse_3_1164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_1165", delete_Data_3_1165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_1166", delete_Found_1166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1167", delete_Key_1167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1168", delete_FoundKey_1168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1169", delete_Data_1169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1170", delete_BtreeIndex_1170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1171", delete_StuckIndex_1171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1172", delete_MergeSuccess_1172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_index_1173", delete_index_1173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_size_1174", delete_size_1174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isLeaf_1175", delete_isLeaf_1175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_nextFree_1176", delete_nextFree_1176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_0_1177", delete_Key_0_1177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_0_1178", delete_KeyCompares_0_1178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_0_1179", delete_KeyCollapse_0_1179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_0_1180", delete_Data_0_1180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1_1181", delete_Key_1_1181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_1_1182", delete_KeyCompares_1_1182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_1_1183", delete_KeyCollapse_1_1183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1_1184", delete_Data_1_1184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_2_1185", delete_Key_2_1185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_2_1186", delete_KeyCompares_2_1186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_2_1187", delete_KeyCollapse_2_1187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_2_1188", delete_Data_2_1188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_3_1189", delete_Key_3_1189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCompares_3_1190", delete_KeyCompares_3_1190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_KeyCollapse_3_1191", delete_KeyCollapse_3_1191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_3_1192", delete_Data_3_1192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Found_1193", delete_Found_1193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Key_1194", delete_Key_1194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_FoundKey_1195", delete_FoundKey_1195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_Data_1196", delete_Data_1196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_BtreeIndex_1197", delete_BtreeIndex_1197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_StuckIndex_1198", delete_StuckIndex_1198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_MergeSuccess_1199", delete_MergeSuccess_1199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childKey_1200", delete_childKey_1200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_leftChild_1201", delete_leftChild_1201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_rightChild_1202", delete_rightChild_1202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_childData_1203", delete_childData_1203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexLeft_1204", delete_indexLeft_1204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_indexRight_1205", delete_indexRight_1205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_midKey_1206", delete_midKey_1206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_success_1207", delete_success_1207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_test_1208", delete_test_1208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_next_1209", delete_next_1209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_root_1210", delete_root_1210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "delete_isFree_1211", delete_isFree_1211);
      $fclose(o);
    end
  endtask
endmodule
