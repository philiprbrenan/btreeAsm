//-----------------------------------------------------------------------------
// Database on a chip test bench
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree;                                                                      // Test bench for database on a chip
  reg                    stop;                                                  // Program has stopped when this goes high
  reg                   clock;                                                  // Clock
  integer                step;                                                  // Step of the simulation
  integer            maxSteps;                                                  // Maximum number of steps to execute
  integer          returnCode;                                                  // Return code
  integer      processCurrent;                                                  // To ensure we get the same results in Java and Verilog we have to run the processes single threaded in a constant order

  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_stop||stuckData_stop||put_stop;                                                             // Or of process stop fields

  initial begin
    returnCode = 0;
    maxSteps = 200000;
    for(step = -1; step < 0 || step < maxSteps && !stop; step = step + 1) begin // Steps below zero are run unconditionally to initialize each process so that Java and Verilog start in sync at step zero

      processCurrent = 0; clock = 0; #1; clock = 1; #1; // process_stuckIsLeaf_0000
      processCurrent = 1; clock = 0; #1; clock = 1; #1; // process_stuckIsFree_0001
      processCurrent = 2; clock = 0; #1; clock = 1; #1; // process_freeNext_0002
      processCurrent = 3; clock = 0; #1; clock = 1; #1; // process_stuckSize_0003
      processCurrent = 4; clock = 0; #1; clock = 1; #1; // process_stuckKeys_0004
      processCurrent = 5; clock = 0; #1; clock = 1; #1; // process_stuckData_0005
      processCurrent = 6; clock = 0; #1; clock = 1; #1; // process_put_0006
      if (step >= 0) chipPrint();                                            // Steps prior to zero are for initialization to make Java and Verilog match
    end
    if (!stop) $finish(1); else $finish(0);                                // Set return code depending on whether the simulation halted
  end
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[32*1];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_7_result_0;
  integer stuckIsLeaf_7_requestedAt;
  integer stuckIsLeaf_7_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_7_returnCode;
  integer stuckIsLeaf_8_requestedAt;
  integer stuckIsLeaf_8_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_8_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  integer stuckIsLeaf_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_7_result_0 <= 0;
      stuckIsLeaf_7_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_7_returnCode <= 0;
      stuckIsLeaf_8_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_8_returnCode <= 0;
      stuckIsLeaf_memory[0] <= 1;
      for(stuckIsLeaf_memory_index = 1; stuckIsLeaf_memory_index < 32; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
    end
    else if (processCurrent == 0) begin
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_7_result_0 <= stuckIsLeaf_memory[put_stuckIsLeaf_7_index_39*1+0];
            stuckIsLeaf_7_finishedAt <= step;
          end
          else if ((stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step)) begin
            stuckIsLeaf_memory[put_stuckIsLeaf_8_index_40*1+0] <= put_stuckIsLeaf_8_value_41;
            stuckIsLeaf_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[32*1];
  integer stuckIsFree_11_requestedAt;
  integer stuckIsFree_11_finishedAt;
  integer stuckIsFree_stuckIsFree_11_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  integer stuckIsFree_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_11_finishedAt <= -1;
      stuckIsFree_stuckIsFree_11_returnCode <= 0;
      for(stuckIsFree_memory_index = 0; stuckIsFree_memory_index < 1; stuckIsFree_memory_index = stuckIsFree_memory_index + 1) stuckIsFree_memory[stuckIsFree_memory_index] <= 0;
      stuckIsFree_memory[1] <= 1;
      stuckIsFree_memory[2] <= 1;
      stuckIsFree_memory[3] <= 1;
      stuckIsFree_memory[4] <= 1;
      stuckIsFree_memory[5] <= 1;
      stuckIsFree_memory[6] <= 1;
      stuckIsFree_memory[7] <= 1;
      stuckIsFree_memory[8] <= 1;
      stuckIsFree_memory[9] <= 1;
      stuckIsFree_memory[10] <= 1;
      stuckIsFree_memory[11] <= 1;
      stuckIsFree_memory[12] <= 1;
      stuckIsFree_memory[13] <= 1;
      stuckIsFree_memory[14] <= 1;
      stuckIsFree_memory[15] <= 1;
      stuckIsFree_memory[16] <= 1;
      stuckIsFree_memory[17] <= 1;
      stuckIsFree_memory[18] <= 1;
      stuckIsFree_memory[19] <= 1;
      stuckIsFree_memory[20] <= 1;
      stuckIsFree_memory[21] <= 1;
      stuckIsFree_memory[22] <= 1;
      stuckIsFree_memory[23] <= 1;
      stuckIsFree_memory[24] <= 1;
      stuckIsFree_memory[25] <= 1;
      stuckIsFree_memory[26] <= 1;
      stuckIsFree_memory[27] <= 1;
      stuckIsFree_memory[28] <= 1;
      stuckIsFree_memory[29] <= 1;
      stuckIsFree_memory[30] <= 1;
      stuckIsFree_memory[31] <= 1;
    end
    else if (processCurrent == 1) begin
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step)) begin
            stuckIsFree_memory[put_stuckIsFree_11_index_197*1+0] <= put_stuckIsFree_11_value_198;
            stuckIsFree_11_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [6-1:0] freeNext_memory[32*1];
  reg [6-1:0] freeNext_freeNext_9_result_0;
  integer freeNext_9_requestedAt;
  integer freeNext_9_finishedAt;
  integer freeNext_freeNext_9_returnCode;
  integer freeNext_10_requestedAt;
  integer freeNext_10_finishedAt;
  integer freeNext_freeNext_10_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  integer freeNext_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_9_result_0 <= 0;
      freeNext_9_finishedAt <= -1;
      freeNext_freeNext_9_returnCode <= 0;
      freeNext_10_finishedAt <= -1;
      freeNext_freeNext_10_returnCode <= 0;
      freeNext_memory[0] <= 1;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 7;
      freeNext_memory[7] <= 8;
      freeNext_memory[8] <= 9;
      freeNext_memory[9] <= 10;
      freeNext_memory[10] <= 11;
      freeNext_memory[11] <= 12;
      freeNext_memory[12] <= 13;
      freeNext_memory[13] <= 14;
      freeNext_memory[14] <= 15;
      freeNext_memory[15] <= 16;
      freeNext_memory[16] <= 17;
      freeNext_memory[17] <= 18;
      freeNext_memory[18] <= 19;
      freeNext_memory[19] <= 20;
      freeNext_memory[20] <= 21;
      freeNext_memory[21] <= 22;
      freeNext_memory[22] <= 23;
      freeNext_memory[23] <= 24;
      freeNext_memory[24] <= 25;
      freeNext_memory[25] <= 26;
      freeNext_memory[26] <= 27;
      freeNext_memory[27] <= 28;
      freeNext_memory[28] <= 29;
      freeNext_memory[29] <= 30;
      freeNext_memory[30] <= 31;
      for(freeNext_memory_index = 31; freeNext_memory_index < 32; freeNext_memory_index = freeNext_memory_index + 1) freeNext_memory[freeNext_memory_index] <= 0;
    end
    else if (processCurrent == 2) begin
      case(freeNext_pc)
        0: begin
          if ((freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step)) begin
            freeNext_freeNext_9_result_0 <= freeNext_memory[put_freeNext_9_index_194*1+0];
            freeNext_9_finishedAt <= step;
          end
          else if ((freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step)) begin
            freeNext_memory[put_freeNext_10_index_195*1+0] <= put_freeNext_10_value_196;
            freeNext_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[32*1];
  reg [3-1:0] stuckSize_stuckSize_5_result_0;
  integer stuckSize_5_requestedAt;
  integer stuckSize_5_finishedAt;
  integer stuckSize_stuckSize_5_returnCode;
  integer stuckSize_6_requestedAt;
  integer stuckSize_6_finishedAt;
  integer stuckSize_stuckSize_6_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  integer stuckSize_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_5_result_0 <= 0;
      stuckSize_5_finishedAt <= -1;
      stuckSize_stuckSize_5_returnCode <= 0;
      stuckSize_6_finishedAt <= -1;
      stuckSize_stuckSize_6_returnCode <= 0;
      for(stuckSize_memory_index = 0; stuckSize_memory_index < 32; stuckSize_memory_index = stuckSize_memory_index + 1) stuckSize_memory[stuckSize_memory_index] <= 0;
    end
    else if (processCurrent == 3) begin
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step)) begin
            stuckSize_stuckSize_5_result_0 <= stuckSize_memory[put_stuckSize_5_index_36*1+0];
            stuckSize_5_finishedAt <= step;
          end
          else if ((stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step)) begin
            stuckSize_memory[put_stuckSize_6_index_37*1+0] <= put_stuckSize_6_value_38;
            stuckSize_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys  process_stuckKeys_0004
  (* ram_style = "block" *)
  reg [8-1:0] stuckKeys_memory[32*4];
  reg [8-1:0] stuckKeys_stuckKeys_1_result_0;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_1;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_2;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_3;
  integer stuckKeys_1_requestedAt;
  integer stuckKeys_1_finishedAt;
  integer stuckKeys_stuckKeys_1_returnCode;
  integer stuckKeys_2_requestedAt;
  integer stuckKeys_2_finishedAt;
  integer stuckKeys_stuckKeys_2_returnCode;
  integer stuckKeys_pc;
  integer stuckKeys_stop;
  integer stuckKeys_returnCode;
  integer stuckKeys_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_pc <= 0;
      stuckKeys_stop <= 0;
      stuckKeys_returnCode <= 0;
      stuckKeys_stuckKeys_1_result_0 <= 0;
      stuckKeys_stuckKeys_1_result_1 <= 0;
      stuckKeys_stuckKeys_1_result_2 <= 0;
      stuckKeys_stuckKeys_1_result_3 <= 0;
      stuckKeys_1_finishedAt <= -1;
      stuckKeys_stuckKeys_1_returnCode <= 0;
      stuckKeys_2_finishedAt <= -1;
      stuckKeys_stuckKeys_2_returnCode <= 0;
      for(stuckKeys_memory_index = 0; stuckKeys_memory_index < 128; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
    end
    else if (processCurrent == 4) begin
      case(stuckKeys_pc)
        0: begin
          if ((stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step)) begin
            stuckKeys_stuckKeys_1_result_0 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+0];
            stuckKeys_stuckKeys_1_result_1 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+1];
            stuckKeys_stuckKeys_1_result_2 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+2];
            stuckKeys_stuckKeys_1_result_3 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+3];
            stuckKeys_1_finishedAt <= step;
          end
          else if ((stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step)) begin
            stuckKeys_memory[put_stuckKeys_2_index_25*4+0] <= put_stuckKeys_2_value_26;
            stuckKeys_memory[put_stuckKeys_2_index_25*4+1] <= put_stuckKeys_2_value_27;
            stuckKeys_memory[put_stuckKeys_2_index_25*4+2] <= put_stuckKeys_2_value_28;
            stuckKeys_memory[put_stuckKeys_2_index_25*4+3] <= put_stuckKeys_2_value_29;
            stuckKeys_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_stop <= 1;
      endcase
    end
  end
  // Process: stuckData  process_stuckData_0005
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_memory[32*4];
  reg [8-1:0] stuckData_stuckData_3_result_0;
  reg [8-1:0] stuckData_stuckData_3_result_1;
  reg [8-1:0] stuckData_stuckData_3_result_2;
  reg [8-1:0] stuckData_stuckData_3_result_3;
  integer stuckData_3_requestedAt;
  integer stuckData_3_finishedAt;
  integer stuckData_stuckData_3_returnCode;
  integer stuckData_4_requestedAt;
  integer stuckData_4_finishedAt;
  integer stuckData_stuckData_4_returnCode;
  integer stuckData_pc;
  integer stuckData_stop;
  integer stuckData_returnCode;
  integer stuckData_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_pc <= 0;
      stuckData_stop <= 0;
      stuckData_returnCode <= 0;
      stuckData_stuckData_3_result_0 <= 0;
      stuckData_stuckData_3_result_1 <= 0;
      stuckData_stuckData_3_result_2 <= 0;
      stuckData_stuckData_3_result_3 <= 0;
      stuckData_3_finishedAt <= -1;
      stuckData_stuckData_3_returnCode <= 0;
      stuckData_4_finishedAt <= -1;
      stuckData_stuckData_4_returnCode <= 0;
      for(stuckData_memory_index = 0; stuckData_memory_index < 128; stuckData_memory_index = stuckData_memory_index + 1) stuckData_memory[stuckData_memory_index] <= 0;
    end
    else if (processCurrent == 5) begin
      case(stuckData_pc)
        0: begin
          if ((stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step)) begin
            stuckData_stuckData_3_result_0 <= stuckData_memory[put_stuckData_3_index_30*4+0];
            stuckData_stuckData_3_result_1 <= stuckData_memory[put_stuckData_3_index_30*4+1];
            stuckData_stuckData_3_result_2 <= stuckData_memory[put_stuckData_3_index_30*4+2];
            stuckData_stuckData_3_result_3 <= stuckData_memory[put_stuckData_3_index_30*4+3];
            stuckData_3_finishedAt <= step;
          end
          else if ((stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step)) begin
            stuckData_memory[put_stuckData_4_index_31*4+0] <= put_stuckData_4_value_32;
            stuckData_memory[put_stuckData_4_index_31*4+1] <= put_stuckData_4_value_33;
            stuckData_memory[put_stuckData_4_index_31*4+2] <= put_stuckData_4_value_34;
            stuckData_memory[put_stuckData_4_index_31*4+3] <= put_stuckData_4_value_35;
            stuckData_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_stop <= 1;
      endcase
    end
  end
  // Process: put  process_put_0006
  reg [8-1:0] put_k_0;
  reg [8-1:0] put_d_1;
  reg [8-1:0] put_i_2;
  reg [1-1:0] put_l_3;
  reg [6-1:0] put_index_4;
  reg [3-1:0] put_size_5;
  reg [1-1:0] put_isLeaf_6;
  reg [6-1:0] put_nextFree_7;
  reg [8-1:0] put_Key_0_8;
  reg [1-1:0] put_KeyCompares_0_9;
  reg [3-1:0] put_KeyCollapse_0_10;
  reg [8-1:0] put_Data_0_11;
  reg [8-1:0] put_Key_1_12;
  reg [1-1:0] put_KeyCompares_1_13;
  reg [3-1:0] put_KeyCollapse_1_14;
  reg [8-1:0] put_Data_1_15;
  reg [8-1:0] put_Key_2_16;
  reg [1-1:0] put_KeyCompares_2_17;
  reg [3-1:0] put_KeyCollapse_2_18;
  reg [8-1:0] put_Data_2_19;
  reg [8-1:0] put_Key_3_20;
  reg [1-1:0] put_KeyCompares_3_21;
  reg [3-1:0] put_KeyCollapse_3_22;
  reg [8-1:0] put_Data_3_23;
  reg [5-1:0] put_stuckKeys_1_index_24;
  reg [5-1:0] put_stuckKeys_2_index_25;
  reg [8-1:0] put_stuckKeys_2_value_26;
  reg [8-1:0] put_stuckKeys_2_value_27;
  reg [8-1:0] put_stuckKeys_2_value_28;
  reg [8-1:0] put_stuckKeys_2_value_29;
  reg [5-1:0] put_stuckData_3_index_30;
  reg [5-1:0] put_stuckData_4_index_31;
  reg [8-1:0] put_stuckData_4_value_32;
  reg [8-1:0] put_stuckData_4_value_33;
  reg [8-1:0] put_stuckData_4_value_34;
  reg [8-1:0] put_stuckData_4_value_35;
  reg [5-1:0] put_stuckSize_5_index_36;
  reg [5-1:0] put_stuckSize_6_index_37;
  reg [3-1:0] put_stuckSize_6_value_38;
  reg [5-1:0] put_stuckIsLeaf_7_index_39;
  reg [5-1:0] put_stuckIsLeaf_8_index_40;
  reg [1-1:0] put_stuckIsLeaf_8_value_41;
  reg [1-1:0] put_Found_42;
  reg [8-1:0] put_Key_43;
  reg [8-1:0] put_FoundKey_44;
  reg [8-1:0] put_Data_45;
  reg [6-1:0] put_BtreeIndex_46;
  reg [3-1:0] put_StuckIndex_47;
  reg [1-1:0] put_MergeSuccess_48;
  reg [6-1:0] put_index_49;
  reg [3-1:0] put_size_50;
  reg [1-1:0] put_isLeaf_51;
  reg [6-1:0] put_nextFree_52;
  reg [8-1:0] put_Key_0_53;
  reg [1-1:0] put_KeyCompares_0_54;
  reg [3-1:0] put_KeyCollapse_0_55;
  reg [8-1:0] put_Data_0_56;
  reg [8-1:0] put_Key_1_57;
  reg [1-1:0] put_KeyCompares_1_58;
  reg [3-1:0] put_KeyCollapse_1_59;
  reg [8-1:0] put_Data_1_60;
  reg [8-1:0] put_Key_2_61;
  reg [1-1:0] put_KeyCompares_2_62;
  reg [3-1:0] put_KeyCollapse_2_63;
  reg [8-1:0] put_Data_2_64;
  reg [8-1:0] put_Key_3_65;
  reg [1-1:0] put_KeyCompares_3_66;
  reg [3-1:0] put_KeyCollapse_3_67;
  reg [8-1:0] put_Data_3_68;
  reg [1-1:0] put_Found_69;
  reg [8-1:0] put_Key_70;
  reg [8-1:0] put_FoundKey_71;
  reg [8-1:0] put_Data_72;
  reg [6-1:0] put_BtreeIndex_73;
  reg [3-1:0] put_StuckIndex_74;
  reg [1-1:0] put_MergeSuccess_75;
  reg [6-1:0] put_index_76;
  reg [3-1:0] put_size_77;
  reg [1-1:0] put_isLeaf_78;
  reg [6-1:0] put_nextFree_79;
  reg [8-1:0] put_Key_0_80;
  reg [1-1:0] put_KeyCompares_0_81;
  reg [3-1:0] put_KeyCollapse_0_82;
  reg [8-1:0] put_Data_0_83;
  reg [8-1:0] put_Key_1_84;
  reg [1-1:0] put_KeyCompares_1_85;
  reg [3-1:0] put_KeyCollapse_1_86;
  reg [8-1:0] put_Data_1_87;
  reg [8-1:0] put_Key_2_88;
  reg [1-1:0] put_KeyCompares_2_89;
  reg [3-1:0] put_KeyCollapse_2_90;
  reg [8-1:0] put_Data_2_91;
  reg [8-1:0] put_Key_3_92;
  reg [1-1:0] put_KeyCompares_3_93;
  reg [3-1:0] put_KeyCollapse_3_94;
  reg [8-1:0] put_Data_3_95;
  reg [1-1:0] put_Found_96;
  reg [8-1:0] put_Key_97;
  reg [8-1:0] put_FoundKey_98;
  reg [8-1:0] put_Data_99;
  reg [6-1:0] put_BtreeIndex_100;
  reg [3-1:0] put_StuckIndex_101;
  reg [1-1:0] put_MergeSuccess_102;
  reg [6-1:0] put_child_103;
  reg [6-1:0] put_parent_104;
  reg [3-1:0] put_childInparent_105;
  reg [1-1:0] put_found_106;
  reg [1-1:0] put_full_107;
  reg [3-1:0] put_i_108;
  reg [1-1:0] put_notFull_109;
  reg [6-1:0] put_index_110;
  reg [3-1:0] put_size_111;
  reg [1-1:0] put_isLeaf_112;
  reg [6-1:0] put_nextFree_113;
  reg [8-1:0] put_Key_0_114;
  reg [1-1:0] put_KeyCompares_0_115;
  reg [3-1:0] put_KeyCollapse_0_116;
  reg [8-1:0] put_Data_0_117;
  reg [8-1:0] put_Key_1_118;
  reg [1-1:0] put_KeyCompares_1_119;
  reg [3-1:0] put_KeyCollapse_1_120;
  reg [8-1:0] put_Data_1_121;
  reg [8-1:0] put_Key_2_122;
  reg [1-1:0] put_KeyCompares_2_123;
  reg [3-1:0] put_KeyCollapse_2_124;
  reg [8-1:0] put_Data_2_125;
  reg [8-1:0] put_Key_3_126;
  reg [1-1:0] put_KeyCompares_3_127;
  reg [3-1:0] put_KeyCollapse_3_128;
  reg [8-1:0] put_Data_3_129;
  reg [1-1:0] put_Found_130;
  reg [8-1:0] put_Key_131;
  reg [8-1:0] put_FoundKey_132;
  reg [8-1:0] put_Data_133;
  reg [6-1:0] put_BtreeIndex_134;
  reg [3-1:0] put_StuckIndex_135;
  reg [1-1:0] put_MergeSuccess_136;
  reg [6-1:0] put_index_137;
  reg [3-1:0] put_size_138;
  reg [1-1:0] put_isLeaf_139;
  reg [6-1:0] put_nextFree_140;
  reg [8-1:0] put_Key_0_141;
  reg [1-1:0] put_KeyCompares_0_142;
  reg [3-1:0] put_KeyCollapse_0_143;
  reg [8-1:0] put_Data_0_144;
  reg [8-1:0] put_Key_1_145;
  reg [1-1:0] put_KeyCompares_1_146;
  reg [3-1:0] put_KeyCollapse_1_147;
  reg [8-1:0] put_Data_1_148;
  reg [8-1:0] put_Key_2_149;
  reg [1-1:0] put_KeyCompares_2_150;
  reg [3-1:0] put_KeyCollapse_2_151;
  reg [8-1:0] put_Data_2_152;
  reg [8-1:0] put_Key_3_153;
  reg [1-1:0] put_KeyCompares_3_154;
  reg [3-1:0] put_KeyCollapse_3_155;
  reg [8-1:0] put_Data_3_156;
  reg [1-1:0] put_Found_157;
  reg [8-1:0] put_Key_158;
  reg [8-1:0] put_FoundKey_159;
  reg [8-1:0] put_Data_160;
  reg [6-1:0] put_BtreeIndex_161;
  reg [3-1:0] put_StuckIndex_162;
  reg [1-1:0] put_MergeSuccess_163;
  reg [6-1:0] put_index_164;
  reg [3-1:0] put_size_165;
  reg [1-1:0] put_isLeaf_166;
  reg [6-1:0] put_nextFree_167;
  reg [8-1:0] put_Key_0_168;
  reg [1-1:0] put_KeyCompares_0_169;
  reg [3-1:0] put_KeyCollapse_0_170;
  reg [8-1:0] put_Data_0_171;
  reg [8-1:0] put_Key_1_172;
  reg [1-1:0] put_KeyCompares_1_173;
  reg [3-1:0] put_KeyCollapse_1_174;
  reg [8-1:0] put_Data_1_175;
  reg [8-1:0] put_Key_2_176;
  reg [1-1:0] put_KeyCompares_2_177;
  reg [3-1:0] put_KeyCollapse_2_178;
  reg [8-1:0] put_Data_2_179;
  reg [8-1:0] put_Key_3_180;
  reg [1-1:0] put_KeyCompares_3_181;
  reg [3-1:0] put_KeyCollapse_3_182;
  reg [8-1:0] put_Data_3_183;
  reg [1-1:0] put_Found_184;
  reg [8-1:0] put_Key_185;
  reg [8-1:0] put_FoundKey_186;
  reg [8-1:0] put_Data_187;
  reg [6-1:0] put_BtreeIndex_188;
  reg [3-1:0] put_StuckIndex_189;
  reg [1-1:0] put_MergeSuccess_190;
  reg [6-1:0] put_indexLeft_191;
  reg [6-1:0] put_indexRight_192;
  reg [8-1:0] put_midKey_193;
  reg [5-1:0] put_freeNext_9_index_194;
  reg [5-1:0] put_freeNext_10_index_195;
  reg [6-1:0] put_freeNext_10_value_196;
  reg [5-1:0] put_stuckIsFree_11_index_197;
  reg [1-1:0] put_stuckIsFree_11_value_198;
  reg [6-1:0] put_root_199;
  reg [6-1:0] put_next_200;
  reg [1-1:0] put_isLeaf_201;
  reg [1-1:0] put_isFree_202;
  reg [6-1:0] put_root_203;
  reg [6-1:0] put_next_204;
  reg [1-1:0] put_isLeaf_205;
  reg [1-1:0] put_isFree_206;
  reg [3-1:0] put_i_207;
  reg [1-1:0] put_notFull_208;
  reg [6-1:0] put_index_209;
  reg [3-1:0] put_size_210;
  reg [1-1:0] put_isLeaf_211;
  reg [6-1:0] put_nextFree_212;
  reg [8-1:0] put_Key_0_213;
  reg [1-1:0] put_KeyCompares_0_214;
  reg [3-1:0] put_KeyCollapse_0_215;
  reg [8-1:0] put_Data_0_216;
  reg [8-1:0] put_Key_1_217;
  reg [1-1:0] put_KeyCompares_1_218;
  reg [3-1:0] put_KeyCollapse_1_219;
  reg [8-1:0] put_Data_1_220;
  reg [8-1:0] put_Key_2_221;
  reg [1-1:0] put_KeyCompares_2_222;
  reg [3-1:0] put_KeyCollapse_2_223;
  reg [8-1:0] put_Data_2_224;
  reg [8-1:0] put_Key_3_225;
  reg [1-1:0] put_KeyCompares_3_226;
  reg [3-1:0] put_KeyCollapse_3_227;
  reg [8-1:0] put_Data_3_228;
  reg [1-1:0] put_Found_229;
  reg [8-1:0] put_Key_230;
  reg [8-1:0] put_FoundKey_231;
  reg [8-1:0] put_Data_232;
  reg [6-1:0] put_BtreeIndex_233;
  reg [3-1:0] put_StuckIndex_234;
  reg [1-1:0] put_MergeSuccess_235;
  reg [6-1:0] put_index_236;
  reg [3-1:0] put_size_237;
  reg [1-1:0] put_isLeaf_238;
  reg [6-1:0] put_nextFree_239;
  reg [8-1:0] put_Key_0_240;
  reg [1-1:0] put_KeyCompares_0_241;
  reg [3-1:0] put_KeyCollapse_0_242;
  reg [8-1:0] put_Data_0_243;
  reg [8-1:0] put_Key_1_244;
  reg [1-1:0] put_KeyCompares_1_245;
  reg [3-1:0] put_KeyCollapse_1_246;
  reg [8-1:0] put_Data_1_247;
  reg [8-1:0] put_Key_2_248;
  reg [1-1:0] put_KeyCompares_2_249;
  reg [3-1:0] put_KeyCollapse_2_250;
  reg [8-1:0] put_Data_2_251;
  reg [8-1:0] put_Key_3_252;
  reg [1-1:0] put_KeyCompares_3_253;
  reg [3-1:0] put_KeyCollapse_3_254;
  reg [8-1:0] put_Data_3_255;
  reg [1-1:0] put_Found_256;
  reg [8-1:0] put_Key_257;
  reg [8-1:0] put_FoundKey_258;
  reg [8-1:0] put_Data_259;
  reg [6-1:0] put_BtreeIndex_260;
  reg [3-1:0] put_StuckIndex_261;
  reg [1-1:0] put_MergeSuccess_262;
  reg [6-1:0] put_index_263;
  reg [3-1:0] put_size_264;
  reg [1-1:0] put_isLeaf_265;
  reg [6-1:0] put_nextFree_266;
  reg [8-1:0] put_Key_0_267;
  reg [1-1:0] put_KeyCompares_0_268;
  reg [3-1:0] put_KeyCollapse_0_269;
  reg [8-1:0] put_Data_0_270;
  reg [8-1:0] put_Key_1_271;
  reg [1-1:0] put_KeyCompares_1_272;
  reg [3-1:0] put_KeyCollapse_1_273;
  reg [8-1:0] put_Data_1_274;
  reg [8-1:0] put_Key_2_275;
  reg [1-1:0] put_KeyCompares_2_276;
  reg [3-1:0] put_KeyCollapse_2_277;
  reg [8-1:0] put_Data_2_278;
  reg [8-1:0] put_Key_3_279;
  reg [1-1:0] put_KeyCompares_3_280;
  reg [3-1:0] put_KeyCollapse_3_281;
  reg [8-1:0] put_Data_3_282;
  reg [1-1:0] put_Found_283;
  reg [8-1:0] put_Key_284;
  reg [8-1:0] put_FoundKey_285;
  reg [8-1:0] put_Data_286;
  reg [6-1:0] put_BtreeIndex_287;
  reg [3-1:0] put_StuckIndex_288;
  reg [1-1:0] put_MergeSuccess_289;
  reg [6-1:0] put_indexLeft_290;
  reg [6-1:0] put_indexRight_291;
  reg [8-1:0] put_midKey_292;
  reg [6-1:0] put_root_293;
  reg [6-1:0] put_next_294;
  reg [1-1:0] put_isLeaf_295;
  reg [1-1:0] put_isFree_296;
  reg [6-1:0] put_root_297;
  reg [6-1:0] put_next_298;
  reg [1-1:0] put_isLeaf_299;
  reg [1-1:0] put_isFree_300;
  reg [6-1:0] put_index_301;
  reg [3-1:0] put_size_302;
  reg [1-1:0] put_isLeaf_303;
  reg [6-1:0] put_nextFree_304;
  reg [8-1:0] put_Key_0_305;
  reg [1-1:0] put_KeyCompares_0_306;
  reg [3-1:0] put_KeyCollapse_0_307;
  reg [8-1:0] put_Data_0_308;
  reg [8-1:0] put_Key_1_309;
  reg [1-1:0] put_KeyCompares_1_310;
  reg [3-1:0] put_KeyCollapse_1_311;
  reg [8-1:0] put_Data_1_312;
  reg [8-1:0] put_Key_2_313;
  reg [1-1:0] put_KeyCompares_2_314;
  reg [3-1:0] put_KeyCollapse_2_315;
  reg [8-1:0] put_Data_2_316;
  reg [8-1:0] put_Key_3_317;
  reg [1-1:0] put_KeyCompares_3_318;
  reg [3-1:0] put_KeyCollapse_3_319;
  reg [8-1:0] put_Data_3_320;
  reg [1-1:0] put_Found_321;
  reg [8-1:0] put_Key_322;
  reg [8-1:0] put_FoundKey_323;
  reg [8-1:0] put_Data_324;
  reg [6-1:0] put_BtreeIndex_325;
  reg [3-1:0] put_StuckIndex_326;
  reg [1-1:0] put_MergeSuccess_327;
  reg [6-1:0] put_index_328;
  reg [3-1:0] put_size_329;
  reg [1-1:0] put_isLeaf_330;
  reg [6-1:0] put_nextFree_331;
  reg [8-1:0] put_Key_0_332;
  reg [1-1:0] put_KeyCompares_0_333;
  reg [3-1:0] put_KeyCollapse_0_334;
  reg [8-1:0] put_Data_0_335;
  reg [8-1:0] put_Key_1_336;
  reg [1-1:0] put_KeyCompares_1_337;
  reg [3-1:0] put_KeyCollapse_1_338;
  reg [8-1:0] put_Data_1_339;
  reg [8-1:0] put_Key_2_340;
  reg [1-1:0] put_KeyCompares_2_341;
  reg [3-1:0] put_KeyCollapse_2_342;
  reg [8-1:0] put_Data_2_343;
  reg [8-1:0] put_Key_3_344;
  reg [1-1:0] put_KeyCompares_3_345;
  reg [3-1:0] put_KeyCollapse_3_346;
  reg [8-1:0] put_Data_3_347;
  reg [1-1:0] put_Found_348;
  reg [8-1:0] put_Key_349;
  reg [8-1:0] put_FoundKey_350;
  reg [8-1:0] put_Data_351;
  reg [6-1:0] put_BtreeIndex_352;
  reg [3-1:0] put_StuckIndex_353;
  reg [1-1:0] put_MergeSuccess_354;
  reg [6-1:0] put_index_355;
  reg [3-1:0] put_size_356;
  reg [1-1:0] put_isLeaf_357;
  reg [6-1:0] put_nextFree_358;
  reg [8-1:0] put_Key_0_359;
  reg [1-1:0] put_KeyCompares_0_360;
  reg [3-1:0] put_KeyCollapse_0_361;
  reg [8-1:0] put_Data_0_362;
  reg [8-1:0] put_Key_1_363;
  reg [1-1:0] put_KeyCompares_1_364;
  reg [3-1:0] put_KeyCollapse_1_365;
  reg [8-1:0] put_Data_1_366;
  reg [8-1:0] put_Key_2_367;
  reg [1-1:0] put_KeyCompares_2_368;
  reg [3-1:0] put_KeyCollapse_2_369;
  reg [8-1:0] put_Data_2_370;
  reg [8-1:0] put_Key_3_371;
  reg [1-1:0] put_KeyCompares_3_372;
  reg [3-1:0] put_KeyCollapse_3_373;
  reg [8-1:0] put_Data_3_374;
  reg [1-1:0] put_Found_375;
  reg [8-1:0] put_Key_376;
  reg [8-1:0] put_FoundKey_377;
  reg [8-1:0] put_Data_378;
  reg [6-1:0] put_BtreeIndex_379;
  reg [3-1:0] put_StuckIndex_380;
  reg [1-1:0] put_MergeSuccess_381;
  reg [6-1:0] put_index_382;
  reg [3-1:0] put_size_383;
  reg [1-1:0] put_isLeaf_384;
  reg [6-1:0] put_nextFree_385;
  reg [8-1:0] put_Key_0_386;
  reg [1-1:0] put_KeyCompares_0_387;
  reg [3-1:0] put_KeyCollapse_0_388;
  reg [8-1:0] put_Data_0_389;
  reg [8-1:0] put_Key_1_390;
  reg [1-1:0] put_KeyCompares_1_391;
  reg [3-1:0] put_KeyCollapse_1_392;
  reg [8-1:0] put_Data_1_393;
  reg [8-1:0] put_Key_2_394;
  reg [1-1:0] put_KeyCompares_2_395;
  reg [3-1:0] put_KeyCollapse_2_396;
  reg [8-1:0] put_Data_2_397;
  reg [8-1:0] put_Key_3_398;
  reg [1-1:0] put_KeyCompares_3_399;
  reg [3-1:0] put_KeyCollapse_3_400;
  reg [8-1:0] put_Data_3_401;
  reg [1-1:0] put_Found_402;
  reg [8-1:0] put_Key_403;
  reg [8-1:0] put_FoundKey_404;
  reg [8-1:0] put_Data_405;
  reg [6-1:0] put_BtreeIndex_406;
  reg [3-1:0] put_StuckIndex_407;
  reg [1-1:0] put_MergeSuccess_408;
  reg [8-1:0] put_childKey_409;
  reg [6-1:0] put_childData_410;
  reg [6-1:0] put_indexLeft_411;
  reg [6-1:0] put_indexRight_412;
  reg [8-1:0] put_midKey_413;
  reg [6-1:0] put_root_414;
  reg [6-1:0] put_next_415;
  reg [1-1:0] put_isLeaf_416;
  reg [1-1:0] put_isFree_417;
  reg [6-1:0] put_index_418;
  reg [3-1:0] put_size_419;
  reg [1-1:0] put_isLeaf_420;
  reg [6-1:0] put_nextFree_421;
  reg [8-1:0] put_Key_0_422;
  reg [1-1:0] put_KeyCompares_0_423;
  reg [3-1:0] put_KeyCollapse_0_424;
  reg [8-1:0] put_Data_0_425;
  reg [8-1:0] put_Key_1_426;
  reg [1-1:0] put_KeyCompares_1_427;
  reg [3-1:0] put_KeyCollapse_1_428;
  reg [8-1:0] put_Data_1_429;
  reg [8-1:0] put_Key_2_430;
  reg [1-1:0] put_KeyCompares_2_431;
  reg [3-1:0] put_KeyCollapse_2_432;
  reg [8-1:0] put_Data_2_433;
  reg [8-1:0] put_Key_3_434;
  reg [1-1:0] put_KeyCompares_3_435;
  reg [3-1:0] put_KeyCollapse_3_436;
  reg [8-1:0] put_Data_3_437;
  reg [1-1:0] put_Found_438;
  reg [8-1:0] put_Key_439;
  reg [8-1:0] put_FoundKey_440;
  reg [8-1:0] put_Data_441;
  reg [6-1:0] put_BtreeIndex_442;
  reg [3-1:0] put_StuckIndex_443;
  reg [1-1:0] put_MergeSuccess_444;
  reg [6-1:0] put_index_445;
  reg [3-1:0] put_size_446;
  reg [1-1:0] put_isLeaf_447;
  reg [6-1:0] put_nextFree_448;
  reg [8-1:0] put_Key_0_449;
  reg [1-1:0] put_KeyCompares_0_450;
  reg [3-1:0] put_KeyCollapse_0_451;
  reg [8-1:0] put_Data_0_452;
  reg [8-1:0] put_Key_1_453;
  reg [1-1:0] put_KeyCompares_1_454;
  reg [3-1:0] put_KeyCollapse_1_455;
  reg [8-1:0] put_Data_1_456;
  reg [8-1:0] put_Key_2_457;
  reg [1-1:0] put_KeyCompares_2_458;
  reg [3-1:0] put_KeyCollapse_2_459;
  reg [8-1:0] put_Data_2_460;
  reg [8-1:0] put_Key_3_461;
  reg [1-1:0] put_KeyCompares_3_462;
  reg [3-1:0] put_KeyCollapse_3_463;
  reg [8-1:0] put_Data_3_464;
  reg [1-1:0] put_Found_465;
  reg [8-1:0] put_Key_466;
  reg [8-1:0] put_FoundKey_467;
  reg [8-1:0] put_Data_468;
  reg [6-1:0] put_BtreeIndex_469;
  reg [3-1:0] put_StuckIndex_470;
  reg [1-1:0] put_MergeSuccess_471;
  reg [6-1:0] put_index_472;
  reg [3-1:0] put_size_473;
  reg [1-1:0] put_isLeaf_474;
  reg [6-1:0] put_nextFree_475;
  reg [8-1:0] put_Key_0_476;
  reg [1-1:0] put_KeyCompares_0_477;
  reg [3-1:0] put_KeyCollapse_0_478;
  reg [8-1:0] put_Data_0_479;
  reg [8-1:0] put_Key_1_480;
  reg [1-1:0] put_KeyCompares_1_481;
  reg [3-1:0] put_KeyCollapse_1_482;
  reg [8-1:0] put_Data_1_483;
  reg [8-1:0] put_Key_2_484;
  reg [1-1:0] put_KeyCompares_2_485;
  reg [3-1:0] put_KeyCollapse_2_486;
  reg [8-1:0] put_Data_2_487;
  reg [8-1:0] put_Key_3_488;
  reg [1-1:0] put_KeyCompares_3_489;
  reg [3-1:0] put_KeyCollapse_3_490;
  reg [8-1:0] put_Data_3_491;
  reg [1-1:0] put_Found_492;
  reg [8-1:0] put_Key_493;
  reg [8-1:0] put_FoundKey_494;
  reg [8-1:0] put_Data_495;
  reg [6-1:0] put_BtreeIndex_496;
  reg [3-1:0] put_StuckIndex_497;
  reg [1-1:0] put_MergeSuccess_498;
  reg [6-1:0] put_childIndex_499;
  reg [6-1:0] put_leftIndex_500;
  reg [8-1:0] put_midKey_501;
  reg [6-1:0] put_root_502;
  reg [6-1:0] put_next_503;
  reg [1-1:0] put_isLeaf_504;
  reg [1-1:0] put_isFree_505;
  reg [3-1:0] put_i_506;
  reg [1-1:0] put_notFull_507;
  reg [6-1:0] put_index_508;
  reg [3-1:0] put_size_509;
  reg [1-1:0] put_isLeaf_510;
  reg [6-1:0] put_nextFree_511;
  reg [8-1:0] put_Key_0_512;
  reg [1-1:0] put_KeyCompares_0_513;
  reg [3-1:0] put_KeyCollapse_0_514;
  reg [8-1:0] put_Data_0_515;
  reg [8-1:0] put_Key_1_516;
  reg [1-1:0] put_KeyCompares_1_517;
  reg [3-1:0] put_KeyCollapse_1_518;
  reg [8-1:0] put_Data_1_519;
  reg [8-1:0] put_Key_2_520;
  reg [1-1:0] put_KeyCompares_2_521;
  reg [3-1:0] put_KeyCollapse_2_522;
  reg [8-1:0] put_Data_2_523;
  reg [8-1:0] put_Key_3_524;
  reg [1-1:0] put_KeyCompares_3_525;
  reg [3-1:0] put_KeyCollapse_3_526;
  reg [8-1:0] put_Data_3_527;
  reg [1-1:0] put_Found_528;
  reg [8-1:0] put_Key_529;
  reg [8-1:0] put_FoundKey_530;
  reg [8-1:0] put_Data_531;
  reg [6-1:0] put_BtreeIndex_532;
  reg [3-1:0] put_StuckIndex_533;
  reg [1-1:0] put_MergeSuccess_534;
  reg [6-1:0] put_index_535;
  reg [3-1:0] put_size_536;
  reg [1-1:0] put_isLeaf_537;
  reg [6-1:0] put_nextFree_538;
  reg [8-1:0] put_Key_0_539;
  reg [1-1:0] put_KeyCompares_0_540;
  reg [3-1:0] put_KeyCollapse_0_541;
  reg [8-1:0] put_Data_0_542;
  reg [8-1:0] put_Key_1_543;
  reg [1-1:0] put_KeyCompares_1_544;
  reg [3-1:0] put_KeyCollapse_1_545;
  reg [8-1:0] put_Data_1_546;
  reg [8-1:0] put_Key_2_547;
  reg [1-1:0] put_KeyCompares_2_548;
  reg [3-1:0] put_KeyCollapse_2_549;
  reg [8-1:0] put_Data_2_550;
  reg [8-1:0] put_Key_3_551;
  reg [1-1:0] put_KeyCompares_3_552;
  reg [3-1:0] put_KeyCollapse_3_553;
  reg [8-1:0] put_Data_3_554;
  reg [1-1:0] put_Found_555;
  reg [8-1:0] put_Key_556;
  reg [8-1:0] put_FoundKey_557;
  reg [8-1:0] put_Data_558;
  reg [6-1:0] put_BtreeIndex_559;
  reg [3-1:0] put_StuckIndex_560;
  reg [1-1:0] put_MergeSuccess_561;
  reg [6-1:0] put_index_562;
  reg [3-1:0] put_size_563;
  reg [1-1:0] put_isLeaf_564;
  reg [6-1:0] put_nextFree_565;
  reg [8-1:0] put_Key_0_566;
  reg [1-1:0] put_KeyCompares_0_567;
  reg [3-1:0] put_KeyCollapse_0_568;
  reg [8-1:0] put_Data_0_569;
  reg [8-1:0] put_Key_1_570;
  reg [1-1:0] put_KeyCompares_1_571;
  reg [3-1:0] put_KeyCollapse_1_572;
  reg [8-1:0] put_Data_1_573;
  reg [8-1:0] put_Key_2_574;
  reg [1-1:0] put_KeyCompares_2_575;
  reg [3-1:0] put_KeyCollapse_2_576;
  reg [8-1:0] put_Data_2_577;
  reg [8-1:0] put_Key_3_578;
  reg [1-1:0] put_KeyCompares_3_579;
  reg [3-1:0] put_KeyCollapse_3_580;
  reg [8-1:0] put_Data_3_581;
  reg [1-1:0] put_Found_582;
  reg [8-1:0] put_Key_583;
  reg [8-1:0] put_FoundKey_584;
  reg [8-1:0] put_Data_585;
  reg [6-1:0] put_BtreeIndex_586;
  reg [3-1:0] put_StuckIndex_587;
  reg [1-1:0] put_MergeSuccess_588;
  reg [6-1:0] put_index_589;
  reg [3-1:0] put_size_590;
  reg [1-1:0] put_isLeaf_591;
  reg [6-1:0] put_nextFree_592;
  reg [8-1:0] put_Key_0_593;
  reg [1-1:0] put_KeyCompares_0_594;
  reg [3-1:0] put_KeyCollapse_0_595;
  reg [8-1:0] put_Data_0_596;
  reg [8-1:0] put_Key_1_597;
  reg [1-1:0] put_KeyCompares_1_598;
  reg [3-1:0] put_KeyCollapse_1_599;
  reg [8-1:0] put_Data_1_600;
  reg [8-1:0] put_Key_2_601;
  reg [1-1:0] put_KeyCompares_2_602;
  reg [3-1:0] put_KeyCollapse_2_603;
  reg [8-1:0] put_Data_2_604;
  reg [8-1:0] put_Key_3_605;
  reg [1-1:0] put_KeyCompares_3_606;
  reg [3-1:0] put_KeyCollapse_3_607;
  reg [8-1:0] put_Data_3_608;
  reg [1-1:0] put_Found_609;
  reg [8-1:0] put_Key_610;
  reg [8-1:0] put_FoundKey_611;
  reg [8-1:0] put_Data_612;
  reg [6-1:0] put_BtreeIndex_613;
  reg [3-1:0] put_StuckIndex_614;
  reg [1-1:0] put_MergeSuccess_615;
  reg [8-1:0] put_childKey_616;
  reg [6-1:0] put_childData_617;
  reg [6-1:0] put_indexLeft_618;
  reg [6-1:0] put_indexRight_619;
  reg [8-1:0] put_midKey_620;
  reg [6-1:0] put_root_621;
  reg [6-1:0] put_next_622;
  reg [1-1:0] put_isLeaf_623;
  reg [1-1:0] put_isFree_624;
  reg [6-1:0] put_index_625;
  reg [3-1:0] put_size_626;
  reg [1-1:0] put_isLeaf_627;
  reg [6-1:0] put_nextFree_628;
  reg [8-1:0] put_Key_0_629;
  reg [1-1:0] put_KeyCompares_0_630;
  reg [3-1:0] put_KeyCollapse_0_631;
  reg [8-1:0] put_Data_0_632;
  reg [8-1:0] put_Key_1_633;
  reg [1-1:0] put_KeyCompares_1_634;
  reg [3-1:0] put_KeyCollapse_1_635;
  reg [8-1:0] put_Data_1_636;
  reg [8-1:0] put_Key_2_637;
  reg [1-1:0] put_KeyCompares_2_638;
  reg [3-1:0] put_KeyCollapse_2_639;
  reg [8-1:0] put_Data_2_640;
  reg [8-1:0] put_Key_3_641;
  reg [1-1:0] put_KeyCompares_3_642;
  reg [3-1:0] put_KeyCollapse_3_643;
  reg [8-1:0] put_Data_3_644;
  reg [1-1:0] put_Found_645;
  reg [8-1:0] put_Key_646;
  reg [8-1:0] put_FoundKey_647;
  reg [8-1:0] put_Data_648;
  reg [6-1:0] put_BtreeIndex_649;
  reg [3-1:0] put_StuckIndex_650;
  reg [1-1:0] put_MergeSuccess_651;
  reg [6-1:0] put_index_652;
  reg [3-1:0] put_size_653;
  reg [1-1:0] put_isLeaf_654;
  reg [6-1:0] put_nextFree_655;
  reg [8-1:0] put_Key_0_656;
  reg [1-1:0] put_KeyCompares_0_657;
  reg [3-1:0] put_KeyCollapse_0_658;
  reg [8-1:0] put_Data_0_659;
  reg [8-1:0] put_Key_1_660;
  reg [1-1:0] put_KeyCompares_1_661;
  reg [3-1:0] put_KeyCollapse_1_662;
  reg [8-1:0] put_Data_1_663;
  reg [8-1:0] put_Key_2_664;
  reg [1-1:0] put_KeyCompares_2_665;
  reg [3-1:0] put_KeyCollapse_2_666;
  reg [8-1:0] put_Data_2_667;
  reg [8-1:0] put_Key_3_668;
  reg [1-1:0] put_KeyCompares_3_669;
  reg [3-1:0] put_KeyCollapse_3_670;
  reg [8-1:0] put_Data_3_671;
  reg [1-1:0] put_Found_672;
  reg [8-1:0] put_Key_673;
  reg [8-1:0] put_FoundKey_674;
  reg [8-1:0] put_Data_675;
  reg [6-1:0] put_BtreeIndex_676;
  reg [3-1:0] put_StuckIndex_677;
  reg [1-1:0] put_MergeSuccess_678;
  reg [6-1:0] put_index_679;
  reg [3-1:0] put_size_680;
  reg [1-1:0] put_isLeaf_681;
  reg [6-1:0] put_nextFree_682;
  reg [8-1:0] put_Key_0_683;
  reg [1-1:0] put_KeyCompares_0_684;
  reg [3-1:0] put_KeyCollapse_0_685;
  reg [8-1:0] put_Data_0_686;
  reg [8-1:0] put_Key_1_687;
  reg [1-1:0] put_KeyCompares_1_688;
  reg [3-1:0] put_KeyCollapse_1_689;
  reg [8-1:0] put_Data_1_690;
  reg [8-1:0] put_Key_2_691;
  reg [1-1:0] put_KeyCompares_2_692;
  reg [3-1:0] put_KeyCollapse_2_693;
  reg [8-1:0] put_Data_2_694;
  reg [8-1:0] put_Key_3_695;
  reg [1-1:0] put_KeyCompares_3_696;
  reg [3-1:0] put_KeyCollapse_3_697;
  reg [8-1:0] put_Data_3_698;
  reg [1-1:0] put_Found_699;
  reg [8-1:0] put_Key_700;
  reg [8-1:0] put_FoundKey_701;
  reg [8-1:0] put_Data_702;
  reg [6-1:0] put_BtreeIndex_703;
  reg [3-1:0] put_StuckIndex_704;
  reg [1-1:0] put_MergeSuccess_705;
  reg [6-1:0] put_index_706;
  reg [3-1:0] put_size_707;
  reg [1-1:0] put_isLeaf_708;
  reg [6-1:0] put_nextFree_709;
  reg [8-1:0] put_Key_0_710;
  reg [1-1:0] put_KeyCompares_0_711;
  reg [3-1:0] put_KeyCollapse_0_712;
  reg [8-1:0] put_Data_0_713;
  reg [8-1:0] put_Key_1_714;
  reg [1-1:0] put_KeyCompares_1_715;
  reg [3-1:0] put_KeyCollapse_1_716;
  reg [8-1:0] put_Data_1_717;
  reg [8-1:0] put_Key_2_718;
  reg [1-1:0] put_KeyCompares_2_719;
  reg [3-1:0] put_KeyCollapse_2_720;
  reg [8-1:0] put_Data_2_721;
  reg [8-1:0] put_Key_3_722;
  reg [1-1:0] put_KeyCompares_3_723;
  reg [3-1:0] put_KeyCollapse_3_724;
  reg [8-1:0] put_Data_3_725;
  reg [1-1:0] put_Found_726;
  reg [8-1:0] put_Key_727;
  reg [8-1:0] put_FoundKey_728;
  reg [8-1:0] put_Data_729;
  reg [6-1:0] put_BtreeIndex_730;
  reg [3-1:0] put_StuckIndex_731;
  reg [1-1:0] put_MergeSuccess_732;
  reg [8-1:0] put_childKey_733;
  reg [6-1:0] put_childData_734;
  reg [6-1:0] put_indexLeft_735;
  reg [6-1:0] put_indexRight_736;
  reg [8-1:0] put_midKey_737;
  reg [6-1:0] put_root_738;
  reg [6-1:0] put_next_739;
  reg [1-1:0] put_isLeaf_740;
  reg [1-1:0] put_isFree_741;
  reg [6-1:0] put_index_742;
  reg [3-1:0] put_size_743;
  reg [1-1:0] put_isLeaf_744;
  reg [6-1:0] put_nextFree_745;
  reg [8-1:0] put_Key_0_746;
  reg [1-1:0] put_KeyCompares_0_747;
  reg [3-1:0] put_KeyCollapse_0_748;
  reg [8-1:0] put_Data_0_749;
  reg [8-1:0] put_Key_1_750;
  reg [1-1:0] put_KeyCompares_1_751;
  reg [3-1:0] put_KeyCollapse_1_752;
  reg [8-1:0] put_Data_1_753;
  reg [8-1:0] put_Key_2_754;
  reg [1-1:0] put_KeyCompares_2_755;
  reg [3-1:0] put_KeyCollapse_2_756;
  reg [8-1:0] put_Data_2_757;
  reg [8-1:0] put_Key_3_758;
  reg [1-1:0] put_KeyCompares_3_759;
  reg [3-1:0] put_KeyCollapse_3_760;
  reg [8-1:0] put_Data_3_761;
  reg [1-1:0] put_Found_762;
  reg [8-1:0] put_Key_763;
  reg [8-1:0] put_FoundKey_764;
  reg [8-1:0] put_Data_765;
  reg [6-1:0] put_BtreeIndex_766;
  reg [3-1:0] put_StuckIndex_767;
  reg [1-1:0] put_MergeSuccess_768;
  reg [6-1:0] put_position_769;
  reg [3-1:0] put_index_770;
  reg [3-1:0] put_index1_771;
  reg [1-1:0] put_within_772;
  reg [1-1:0] put_isLeaf_773;
  reg [6-1:0] put_index_774;
  reg [3-1:0] put_size_775;
  reg [1-1:0] put_isLeaf_776;
  reg [6-1:0] put_nextFree_777;
  reg [8-1:0] put_Key_0_778;
  reg [1-1:0] put_KeyCompares_0_779;
  reg [3-1:0] put_KeyCollapse_0_780;
  reg [8-1:0] put_Data_0_781;
  reg [8-1:0] put_Key_1_782;
  reg [1-1:0] put_KeyCompares_1_783;
  reg [3-1:0] put_KeyCollapse_1_784;
  reg [8-1:0] put_Data_1_785;
  reg [8-1:0] put_Key_2_786;
  reg [1-1:0] put_KeyCompares_2_787;
  reg [3-1:0] put_KeyCollapse_2_788;
  reg [8-1:0] put_Data_2_789;
  reg [8-1:0] put_Key_3_790;
  reg [1-1:0] put_KeyCompares_3_791;
  reg [3-1:0] put_KeyCollapse_3_792;
  reg [8-1:0] put_Data_3_793;
  reg [1-1:0] put_Found_794;
  reg [8-1:0] put_Key_795;
  reg [8-1:0] put_FoundKey_796;
  reg [8-1:0] put_Data_797;
  reg [6-1:0] put_BtreeIndex_798;
  reg [3-1:0] put_StuckIndex_799;
  reg [1-1:0] put_MergeSuccess_800;
  reg [6-1:0] put_index_801;
  reg [3-1:0] put_size_802;
  reg [1-1:0] put_isLeaf_803;
  reg [6-1:0] put_nextFree_804;
  reg [8-1:0] put_Key_0_805;
  reg [1-1:0] put_KeyCompares_0_806;
  reg [3-1:0] put_KeyCollapse_0_807;
  reg [8-1:0] put_Data_0_808;
  reg [8-1:0] put_Key_1_809;
  reg [1-1:0] put_KeyCompares_1_810;
  reg [3-1:0] put_KeyCollapse_1_811;
  reg [8-1:0] put_Data_1_812;
  reg [8-1:0] put_Key_2_813;
  reg [1-1:0] put_KeyCompares_2_814;
  reg [3-1:0] put_KeyCollapse_2_815;
  reg [8-1:0] put_Data_2_816;
  reg [8-1:0] put_Key_3_817;
  reg [1-1:0] put_KeyCompares_3_818;
  reg [3-1:0] put_KeyCollapse_3_819;
  reg [8-1:0] put_Data_3_820;
  reg [1-1:0] put_Found_821;
  reg [8-1:0] put_Key_822;
  reg [8-1:0] put_FoundKey_823;
  reg [8-1:0] put_Data_824;
  reg [6-1:0] put_BtreeIndex_825;
  reg [3-1:0] put_StuckIndex_826;
  reg [1-1:0] put_MergeSuccess_827;
  reg [6-1:0] put_index_828;
  reg [3-1:0] put_size_829;
  reg [1-1:0] put_isLeaf_830;
  reg [6-1:0] put_nextFree_831;
  reg [8-1:0] put_Key_0_832;
  reg [1-1:0] put_KeyCompares_0_833;
  reg [3-1:0] put_KeyCollapse_0_834;
  reg [8-1:0] put_Data_0_835;
  reg [8-1:0] put_Key_1_836;
  reg [1-1:0] put_KeyCompares_1_837;
  reg [3-1:0] put_KeyCollapse_1_838;
  reg [8-1:0] put_Data_1_839;
  reg [8-1:0] put_Key_2_840;
  reg [1-1:0] put_KeyCompares_2_841;
  reg [3-1:0] put_KeyCollapse_2_842;
  reg [8-1:0] put_Data_2_843;
  reg [8-1:0] put_Key_3_844;
  reg [1-1:0] put_KeyCompares_3_845;
  reg [3-1:0] put_KeyCollapse_3_846;
  reg [8-1:0] put_Data_3_847;
  reg [1-1:0] put_Found_848;
  reg [8-1:0] put_Key_849;
  reg [8-1:0] put_FoundKey_850;
  reg [8-1:0] put_Data_851;
  reg [6-1:0] put_BtreeIndex_852;
  reg [3-1:0] put_StuckIndex_853;
  reg [1-1:0] put_MergeSuccess_854;
  reg [8-1:0] put_childKey_855;
  reg [6-1:0] put_childData_856;
  reg [6-1:0] put_indexLeft_857;
  reg [6-1:0] put_indexRight_858;
  reg [8-1:0] put_midKey_859;
  reg [1-1:0] put_success_860;
  reg [1-1:0] put_test_861;
  reg [6-1:0] put_next_862;
  reg [6-1:0] put_root_863;
  reg [1-1:0] put_isFree_864;
  reg [6-1:0] put_next_865;
  reg [6-1:0] put_root_866;
  reg [1-1:0] put_isFree_867;
  reg [6-1:0] put_index_868;
  reg [3-1:0] put_size_869;
  reg [1-1:0] put_isLeaf_870;
  reg [6-1:0] put_nextFree_871;
  reg [8-1:0] put_Key_0_872;
  reg [1-1:0] put_KeyCompares_0_873;
  reg [3-1:0] put_KeyCollapse_0_874;
  reg [8-1:0] put_Data_0_875;
  reg [8-1:0] put_Key_1_876;
  reg [1-1:0] put_KeyCompares_1_877;
  reg [3-1:0] put_KeyCollapse_1_878;
  reg [8-1:0] put_Data_1_879;
  reg [8-1:0] put_Key_2_880;
  reg [1-1:0] put_KeyCompares_2_881;
  reg [3-1:0] put_KeyCollapse_2_882;
  reg [8-1:0] put_Data_2_883;
  reg [8-1:0] put_Key_3_884;
  reg [1-1:0] put_KeyCompares_3_885;
  reg [3-1:0] put_KeyCollapse_3_886;
  reg [8-1:0] put_Data_3_887;
  reg [1-1:0] put_Found_888;
  reg [8-1:0] put_Key_889;
  reg [8-1:0] put_FoundKey_890;
  reg [8-1:0] put_Data_891;
  reg [6-1:0] put_BtreeIndex_892;
  reg [3-1:0] put_StuckIndex_893;
  reg [1-1:0] put_MergeSuccess_894;
  reg [6-1:0] put_index_895;
  reg [3-1:0] put_size_896;
  reg [1-1:0] put_isLeaf_897;
  reg [6-1:0] put_nextFree_898;
  reg [8-1:0] put_Key_0_899;
  reg [1-1:0] put_KeyCompares_0_900;
  reg [3-1:0] put_KeyCollapse_0_901;
  reg [8-1:0] put_Data_0_902;
  reg [8-1:0] put_Key_1_903;
  reg [1-1:0] put_KeyCompares_1_904;
  reg [3-1:0] put_KeyCollapse_1_905;
  reg [8-1:0] put_Data_1_906;
  reg [8-1:0] put_Key_2_907;
  reg [1-1:0] put_KeyCompares_2_908;
  reg [3-1:0] put_KeyCollapse_2_909;
  reg [8-1:0] put_Data_2_910;
  reg [8-1:0] put_Key_3_911;
  reg [1-1:0] put_KeyCompares_3_912;
  reg [3-1:0] put_KeyCollapse_3_913;
  reg [8-1:0] put_Data_3_914;
  reg [1-1:0] put_Found_915;
  reg [8-1:0] put_Key_916;
  reg [8-1:0] put_FoundKey_917;
  reg [8-1:0] put_Data_918;
  reg [6-1:0] put_BtreeIndex_919;
  reg [3-1:0] put_StuckIndex_920;
  reg [1-1:0] put_MergeSuccess_921;
  reg [6-1:0] put_index_922;
  reg [3-1:0] put_size_923;
  reg [1-1:0] put_isLeaf_924;
  reg [6-1:0] put_nextFree_925;
  reg [8-1:0] put_Key_0_926;
  reg [1-1:0] put_KeyCompares_0_927;
  reg [3-1:0] put_KeyCollapse_0_928;
  reg [8-1:0] put_Data_0_929;
  reg [8-1:0] put_Key_1_930;
  reg [1-1:0] put_KeyCompares_1_931;
  reg [3-1:0] put_KeyCollapse_1_932;
  reg [8-1:0] put_Data_1_933;
  reg [8-1:0] put_Key_2_934;
  reg [1-1:0] put_KeyCompares_2_935;
  reg [3-1:0] put_KeyCollapse_2_936;
  reg [8-1:0] put_Data_2_937;
  reg [8-1:0] put_Key_3_938;
  reg [1-1:0] put_KeyCompares_3_939;
  reg [3-1:0] put_KeyCollapse_3_940;
  reg [8-1:0] put_Data_3_941;
  reg [1-1:0] put_Found_942;
  reg [8-1:0] put_Key_943;
  reg [8-1:0] put_FoundKey_944;
  reg [8-1:0] put_Data_945;
  reg [6-1:0] put_BtreeIndex_946;
  reg [3-1:0] put_StuckIndex_947;
  reg [1-1:0] put_MergeSuccess_948;
  reg [8-1:0] put_childKey_949;
  reg [3-1:0] put_leftChild_950;
  reg [3-1:0] put_rightChild_951;
  reg [6-1:0] put_childData_952;
  reg [6-1:0] put_indexLeft_953;
  reg [6-1:0] put_indexRight_954;
  reg [8-1:0] put_midKey_955;
  reg [1-1:0] put_success_956;
  reg [1-1:0] put_test_957;
  reg [6-1:0] put_next_958;
  reg [6-1:0] put_root_959;
  reg [1-1:0] put_isFree_960;
  reg [6-1:0] put_next_961;
  reg [6-1:0] put_root_962;
  reg [1-1:0] put_isFree_963;
  reg [6-1:0] put_index_964;
  reg [3-1:0] put_size_965;
  reg [1-1:0] put_isLeaf_966;
  reg [6-1:0] put_nextFree_967;
  reg [8-1:0] put_Key_0_968;
  reg [1-1:0] put_KeyCompares_0_969;
  reg [3-1:0] put_KeyCollapse_0_970;
  reg [8-1:0] put_Data_0_971;
  reg [8-1:0] put_Key_1_972;
  reg [1-1:0] put_KeyCompares_1_973;
  reg [3-1:0] put_KeyCollapse_1_974;
  reg [8-1:0] put_Data_1_975;
  reg [8-1:0] put_Key_2_976;
  reg [1-1:0] put_KeyCompares_2_977;
  reg [3-1:0] put_KeyCollapse_2_978;
  reg [8-1:0] put_Data_2_979;
  reg [8-1:0] put_Key_3_980;
  reg [1-1:0] put_KeyCompares_3_981;
  reg [3-1:0] put_KeyCollapse_3_982;
  reg [8-1:0] put_Data_3_983;
  reg [1-1:0] put_Found_984;
  reg [8-1:0] put_Key_985;
  reg [8-1:0] put_FoundKey_986;
  reg [8-1:0] put_Data_987;
  reg [6-1:0] put_BtreeIndex_988;
  reg [3-1:0] put_StuckIndex_989;
  reg [1-1:0] put_MergeSuccess_990;
  reg [6-1:0] put_index_991;
  reg [3-1:0] put_size_992;
  reg [1-1:0] put_isLeaf_993;
  reg [6-1:0] put_nextFree_994;
  reg [8-1:0] put_Key_0_995;
  reg [1-1:0] put_KeyCompares_0_996;
  reg [3-1:0] put_KeyCollapse_0_997;
  reg [8-1:0] put_Data_0_998;
  reg [8-1:0] put_Key_1_999;
  reg [1-1:0] put_KeyCompares_1_1000;
  reg [3-1:0] put_KeyCollapse_1_1001;
  reg [8-1:0] put_Data_1_1002;
  reg [8-1:0] put_Key_2_1003;
  reg [1-1:0] put_KeyCompares_2_1004;
  reg [3-1:0] put_KeyCollapse_2_1005;
  reg [8-1:0] put_Data_2_1006;
  reg [8-1:0] put_Key_3_1007;
  reg [1-1:0] put_KeyCompares_3_1008;
  reg [3-1:0] put_KeyCollapse_3_1009;
  reg [8-1:0] put_Data_3_1010;
  reg [1-1:0] put_Found_1011;
  reg [8-1:0] put_Key_1012;
  reg [8-1:0] put_FoundKey_1013;
  reg [8-1:0] put_Data_1014;
  reg [6-1:0] put_BtreeIndex_1015;
  reg [3-1:0] put_StuckIndex_1016;
  reg [1-1:0] put_MergeSuccess_1017;
  reg [8-1:0] put_childKey_1018;
  reg [3-1:0] put_size_1019;
  reg [6-1:0] put_childData_1020;
  reg [6-1:0] put_indexLeft_1021;
  reg [6-1:0] put_indexRight_1022;
  reg [8-1:0] put_midKey_1023;
  reg [1-1:0] put_success_1024;
  reg [1-1:0] put_test_1025;
  reg [6-1:0] put_next_1026;
  reg [6-1:0] put_root_1027;
  reg [1-1:0] put_isFree_1028;
  reg [6-1:0] put_index_1029;
  reg [3-1:0] put_size_1030;
  reg [1-1:0] put_isLeaf_1031;
  reg [6-1:0] put_nextFree_1032;
  reg [8-1:0] put_Key_0_1033;
  reg [1-1:0] put_KeyCompares_0_1034;
  reg [3-1:0] put_KeyCollapse_0_1035;
  reg [8-1:0] put_Data_0_1036;
  reg [8-1:0] put_Key_1_1037;
  reg [1-1:0] put_KeyCompares_1_1038;
  reg [3-1:0] put_KeyCollapse_1_1039;
  reg [8-1:0] put_Data_1_1040;
  reg [8-1:0] put_Key_2_1041;
  reg [1-1:0] put_KeyCompares_2_1042;
  reg [3-1:0] put_KeyCollapse_2_1043;
  reg [8-1:0] put_Data_2_1044;
  reg [8-1:0] put_Key_3_1045;
  reg [1-1:0] put_KeyCompares_3_1046;
  reg [3-1:0] put_KeyCollapse_3_1047;
  reg [8-1:0] put_Data_3_1048;
  reg [1-1:0] put_Found_1049;
  reg [8-1:0] put_Key_1050;
  reg [8-1:0] put_FoundKey_1051;
  reg [8-1:0] put_Data_1052;
  reg [6-1:0] put_BtreeIndex_1053;
  reg [3-1:0] put_StuckIndex_1054;
  reg [1-1:0] put_MergeSuccess_1055;
  reg [6-1:0] put_index_1056;
  reg [3-1:0] put_size_1057;
  reg [1-1:0] put_isLeaf_1058;
  reg [6-1:0] put_nextFree_1059;
  reg [8-1:0] put_Key_0_1060;
  reg [1-1:0] put_KeyCompares_0_1061;
  reg [3-1:0] put_KeyCollapse_0_1062;
  reg [8-1:0] put_Data_0_1063;
  reg [8-1:0] put_Key_1_1064;
  reg [1-1:0] put_KeyCompares_1_1065;
  reg [3-1:0] put_KeyCollapse_1_1066;
  reg [8-1:0] put_Data_1_1067;
  reg [8-1:0] put_Key_2_1068;
  reg [1-1:0] put_KeyCompares_2_1069;
  reg [3-1:0] put_KeyCollapse_2_1070;
  reg [8-1:0] put_Data_2_1071;
  reg [8-1:0] put_Key_3_1072;
  reg [1-1:0] put_KeyCompares_3_1073;
  reg [3-1:0] put_KeyCollapse_3_1074;
  reg [8-1:0] put_Data_3_1075;
  reg [1-1:0] put_Found_1076;
  reg [8-1:0] put_Key_1077;
  reg [8-1:0] put_FoundKey_1078;
  reg [8-1:0] put_Data_1079;
  reg [6-1:0] put_BtreeIndex_1080;
  reg [3-1:0] put_StuckIndex_1081;
  reg [1-1:0] put_MergeSuccess_1082;
  reg [8-1:0] put_childKey_1083;
  reg [3-1:0] put_size_1084;
  reg [6-1:0] put_childData_1085;
  reg [6-1:0] put_indexLeft_1086;
  reg [6-1:0] put_indexRight_1087;
  reg [8-1:0] put_midKey_1088;
  reg [1-1:0] put_success_1089;
  reg [1-1:0] put_test_1090;
  reg [6-1:0] put_next_1091;
  reg [6-1:0] put_root_1092;
  reg [1-1:0] put_isFree_1093;
  reg [6-1:0] put_index_1094;
  reg [3-1:0] put_size_1095;
  reg [1-1:0] put_isLeaf_1096;
  reg [6-1:0] put_nextFree_1097;
  reg [8-1:0] put_Key_0_1098;
  reg [1-1:0] put_KeyCompares_0_1099;
  reg [3-1:0] put_KeyCollapse_0_1100;
  reg [8-1:0] put_Data_0_1101;
  reg [8-1:0] put_Key_1_1102;
  reg [1-1:0] put_KeyCompares_1_1103;
  reg [3-1:0] put_KeyCollapse_1_1104;
  reg [8-1:0] put_Data_1_1105;
  reg [8-1:0] put_Key_2_1106;
  reg [1-1:0] put_KeyCompares_2_1107;
  reg [3-1:0] put_KeyCollapse_2_1108;
  reg [8-1:0] put_Data_2_1109;
  reg [8-1:0] put_Key_3_1110;
  reg [1-1:0] put_KeyCompares_3_1111;
  reg [3-1:0] put_KeyCollapse_3_1112;
  reg [8-1:0] put_Data_3_1113;
  reg [1-1:0] put_Found_1114;
  reg [8-1:0] put_Key_1115;
  reg [8-1:0] put_FoundKey_1116;
  reg [8-1:0] put_Data_1117;
  reg [6-1:0] put_BtreeIndex_1118;
  reg [3-1:0] put_StuckIndex_1119;
  reg [1-1:0] put_MergeSuccess_1120;
  reg [6-1:0] put_index_1121;
  reg [3-1:0] put_size_1122;
  reg [1-1:0] put_isLeaf_1123;
  reg [6-1:0] put_nextFree_1124;
  reg [8-1:0] put_Key_0_1125;
  reg [1-1:0] put_KeyCompares_0_1126;
  reg [3-1:0] put_KeyCollapse_0_1127;
  reg [8-1:0] put_Data_0_1128;
  reg [8-1:0] put_Key_1_1129;
  reg [1-1:0] put_KeyCompares_1_1130;
  reg [3-1:0] put_KeyCollapse_1_1131;
  reg [8-1:0] put_Data_1_1132;
  reg [8-1:0] put_Key_2_1133;
  reg [1-1:0] put_KeyCompares_2_1134;
  reg [3-1:0] put_KeyCollapse_2_1135;
  reg [8-1:0] put_Data_2_1136;
  reg [8-1:0] put_Key_3_1137;
  reg [1-1:0] put_KeyCompares_3_1138;
  reg [3-1:0] put_KeyCollapse_3_1139;
  reg [8-1:0] put_Data_3_1140;
  reg [1-1:0] put_Found_1141;
  reg [8-1:0] put_Key_1142;
  reg [8-1:0] put_FoundKey_1143;
  reg [8-1:0] put_Data_1144;
  reg [6-1:0] put_BtreeIndex_1145;
  reg [3-1:0] put_StuckIndex_1146;
  reg [1-1:0] put_MergeSuccess_1147;
  reg [8-1:0] put_childKey_1148;
  reg [6-1:0] put_childData_1149;
  reg [6-1:0] put_indexLeft_1150;
  reg [6-1:0] put_indexRight_1151;
  reg [8-1:0] put_midKey_1152;
  reg [1-1:0] put_success_1153;
  reg [1-1:0] put_test_1154;
  reg [6-1:0] put_next_1155;
  reg [6-1:0] put_root_1156;
  reg [1-1:0] put_isFree_1157;
  reg [6-1:0] put_index_1158;
  reg [3-1:0] put_size_1159;
  reg [1-1:0] put_isLeaf_1160;
  reg [6-1:0] put_nextFree_1161;
  reg [8-1:0] put_Key_0_1162;
  reg [1-1:0] put_KeyCompares_0_1163;
  reg [3-1:0] put_KeyCollapse_0_1164;
  reg [8-1:0] put_Data_0_1165;
  reg [8-1:0] put_Key_1_1166;
  reg [1-1:0] put_KeyCompares_1_1167;
  reg [3-1:0] put_KeyCollapse_1_1168;
  reg [8-1:0] put_Data_1_1169;
  reg [8-1:0] put_Key_2_1170;
  reg [1-1:0] put_KeyCompares_2_1171;
  reg [3-1:0] put_KeyCollapse_2_1172;
  reg [8-1:0] put_Data_2_1173;
  reg [8-1:0] put_Key_3_1174;
  reg [1-1:0] put_KeyCompares_3_1175;
  reg [3-1:0] put_KeyCollapse_3_1176;
  reg [8-1:0] put_Data_3_1177;
  reg [1-1:0] put_Found_1178;
  reg [8-1:0] put_Key_1179;
  reg [8-1:0] put_FoundKey_1180;
  reg [8-1:0] put_Data_1181;
  reg [6-1:0] put_BtreeIndex_1182;
  reg [3-1:0] put_StuckIndex_1183;
  reg [1-1:0] put_MergeSuccess_1184;
  reg [6-1:0] put_index_1185;
  reg [3-1:0] put_size_1186;
  reg [1-1:0] put_isLeaf_1187;
  reg [6-1:0] put_nextFree_1188;
  reg [8-1:0] put_Key_0_1189;
  reg [1-1:0] put_KeyCompares_0_1190;
  reg [3-1:0] put_KeyCollapse_0_1191;
  reg [8-1:0] put_Data_0_1192;
  reg [8-1:0] put_Key_1_1193;
  reg [1-1:0] put_KeyCompares_1_1194;
  reg [3-1:0] put_KeyCollapse_1_1195;
  reg [8-1:0] put_Data_1_1196;
  reg [8-1:0] put_Key_2_1197;
  reg [1-1:0] put_KeyCompares_2_1198;
  reg [3-1:0] put_KeyCollapse_2_1199;
  reg [8-1:0] put_Data_2_1200;
  reg [8-1:0] put_Key_3_1201;
  reg [1-1:0] put_KeyCompares_3_1202;
  reg [3-1:0] put_KeyCollapse_3_1203;
  reg [8-1:0] put_Data_3_1204;
  reg [1-1:0] put_Found_1205;
  reg [8-1:0] put_Key_1206;
  reg [8-1:0] put_FoundKey_1207;
  reg [8-1:0] put_Data_1208;
  reg [6-1:0] put_BtreeIndex_1209;
  reg [3-1:0] put_StuckIndex_1210;
  reg [1-1:0] put_MergeSuccess_1211;
  reg [8-1:0] put_childKey_1212;
  reg [3-1:0] put_leftChild_1213;
  reg [3-1:0] put_rightChild_1214;
  reg [6-1:0] put_childData_1215;
  reg [6-1:0] put_indexLeft_1216;
  reg [6-1:0] put_indexRight_1217;
  reg [8-1:0] put_midKey_1218;
  reg [1-1:0] put_success_1219;
  reg [1-1:0] put_test_1220;
  reg [6-1:0] put_next_1221;
  reg [6-1:0] put_root_1222;
  reg [1-1:0] put_isFree_1223;
  reg [6-1:0] put_index_1224;
  reg [3-1:0] put_size_1225;
  reg [1-1:0] put_isLeaf_1226;
  reg [6-1:0] put_nextFree_1227;
  reg [8-1:0] put_Key_0_1228;
  reg [1-1:0] put_KeyCompares_0_1229;
  reg [3-1:0] put_KeyCollapse_0_1230;
  reg [8-1:0] put_Data_0_1231;
  reg [8-1:0] put_Key_1_1232;
  reg [1-1:0] put_KeyCompares_1_1233;
  reg [3-1:0] put_KeyCollapse_1_1234;
  reg [8-1:0] put_Data_1_1235;
  reg [8-1:0] put_Key_2_1236;
  reg [1-1:0] put_KeyCompares_2_1237;
  reg [3-1:0] put_KeyCollapse_2_1238;
  reg [8-1:0] put_Data_2_1239;
  reg [8-1:0] put_Key_3_1240;
  reg [1-1:0] put_KeyCompares_3_1241;
  reg [3-1:0] put_KeyCollapse_3_1242;
  reg [8-1:0] put_Data_3_1243;
  reg [1-1:0] put_Found_1244;
  reg [8-1:0] put_Key_1245;
  reg [8-1:0] put_FoundKey_1246;
  reg [8-1:0] put_Data_1247;
  reg [6-1:0] put_BtreeIndex_1248;
  reg [3-1:0] put_StuckIndex_1249;
  reg [1-1:0] put_MergeSuccess_1250;
  reg [6-1:0] put_index_1251;
  reg [3-1:0] put_size_1252;
  reg [1-1:0] put_isLeaf_1253;
  reg [6-1:0] put_nextFree_1254;
  reg [8-1:0] put_Key_0_1255;
  reg [1-1:0] put_KeyCompares_0_1256;
  reg [3-1:0] put_KeyCollapse_0_1257;
  reg [8-1:0] put_Data_0_1258;
  reg [8-1:0] put_Key_1_1259;
  reg [1-1:0] put_KeyCompares_1_1260;
  reg [3-1:0] put_KeyCollapse_1_1261;
  reg [8-1:0] put_Data_1_1262;
  reg [8-1:0] put_Key_2_1263;
  reg [1-1:0] put_KeyCompares_2_1264;
  reg [3-1:0] put_KeyCollapse_2_1265;
  reg [8-1:0] put_Data_2_1266;
  reg [8-1:0] put_Key_3_1267;
  reg [1-1:0] put_KeyCompares_3_1268;
  reg [3-1:0] put_KeyCollapse_3_1269;
  reg [8-1:0] put_Data_3_1270;
  reg [1-1:0] put_Found_1271;
  reg [8-1:0] put_Key_1272;
  reg [8-1:0] put_FoundKey_1273;
  reg [8-1:0] put_Data_1274;
  reg [6-1:0] put_BtreeIndex_1275;
  reg [3-1:0] put_StuckIndex_1276;
  reg [1-1:0] put_MergeSuccess_1277;
  reg [8-1:0] put_childKey_1278;
  reg [6-1:0] put_childData_1279;
  reg [6-1:0] put_indexLeft_1280;
  reg [6-1:0] put_indexRight_1281;
  reg [8-1:0] put_midKey_1282;
  reg [1-1:0] put_success_1283;
  reg [1-1:0] put_test_1284;
  reg [6-1:0] put_next_1285;
  reg [6-1:0] put_root_1286;
  reg [1-1:0] put_isFree_1287;
  reg [6-1:0] put_index_1288;
  reg [3-1:0] put_size_1289;
  reg [1-1:0] put_isLeaf_1290;
  reg [6-1:0] put_nextFree_1291;
  reg [8-1:0] put_Key_0_1292;
  reg [1-1:0] put_KeyCompares_0_1293;
  reg [3-1:0] put_KeyCollapse_0_1294;
  reg [8-1:0] put_Data_0_1295;
  reg [8-1:0] put_Key_1_1296;
  reg [1-1:0] put_KeyCompares_1_1297;
  reg [3-1:0] put_KeyCollapse_1_1298;
  reg [8-1:0] put_Data_1_1299;
  reg [8-1:0] put_Key_2_1300;
  reg [1-1:0] put_KeyCompares_2_1301;
  reg [3-1:0] put_KeyCollapse_2_1302;
  reg [8-1:0] put_Data_2_1303;
  reg [8-1:0] put_Key_3_1304;
  reg [1-1:0] put_KeyCompares_3_1305;
  reg [3-1:0] put_KeyCollapse_3_1306;
  reg [8-1:0] put_Data_3_1307;
  reg [1-1:0] put_Found_1308;
  reg [8-1:0] put_Key_1309;
  reg [8-1:0] put_FoundKey_1310;
  reg [8-1:0] put_Data_1311;
  reg [6-1:0] put_BtreeIndex_1312;
  reg [3-1:0] put_StuckIndex_1313;
  reg [1-1:0] put_MergeSuccess_1314;
  reg [6-1:0] put_index_1315;
  reg [3-1:0] put_size_1316;
  reg [1-1:0] put_isLeaf_1317;
  reg [6-1:0] put_nextFree_1318;
  reg [8-1:0] put_Key_0_1319;
  reg [1-1:0] put_KeyCompares_0_1320;
  reg [3-1:0] put_KeyCollapse_0_1321;
  reg [8-1:0] put_Data_0_1322;
  reg [8-1:0] put_Key_1_1323;
  reg [1-1:0] put_KeyCompares_1_1324;
  reg [3-1:0] put_KeyCollapse_1_1325;
  reg [8-1:0] put_Data_1_1326;
  reg [8-1:0] put_Key_2_1327;
  reg [1-1:0] put_KeyCompares_2_1328;
  reg [3-1:0] put_KeyCollapse_2_1329;
  reg [8-1:0] put_Data_2_1330;
  reg [8-1:0] put_Key_3_1331;
  reg [1-1:0] put_KeyCompares_3_1332;
  reg [3-1:0] put_KeyCollapse_3_1333;
  reg [8-1:0] put_Data_3_1334;
  reg [1-1:0] put_Found_1335;
  reg [8-1:0] put_Key_1336;
  reg [8-1:0] put_FoundKey_1337;
  reg [8-1:0] put_Data_1338;
  reg [6-1:0] put_BtreeIndex_1339;
  reg [3-1:0] put_StuckIndex_1340;
  reg [1-1:0] put_MergeSuccess_1341;
  reg [8-1:0] put_childKey_1342;
  reg [3-1:0] put_leftChild_1343;
  reg [3-1:0] put_rightChild_1344;
  reg [6-1:0] put_childData_1345;
  reg [6-1:0] put_indexLeft_1346;
  reg [6-1:0] put_indexRight_1347;
  reg [8-1:0] put_midKey_1348;
  reg [1-1:0] put_success_1349;
  reg [1-1:0] put_test_1350;
  reg [6-1:0] put_next_1351;
  reg [6-1:0] put_root_1352;
  reg [1-1:0] put_isFree_1353;
  reg [6-1:0] put_index_1354;
  reg [3-1:0] put_size_1355;
  reg [1-1:0] put_isLeaf_1356;
  reg [6-1:0] put_nextFree_1357;
  reg [8-1:0] put_Key_0_1358;
  reg [1-1:0] put_KeyCompares_0_1359;
  reg [3-1:0] put_KeyCollapse_0_1360;
  reg [8-1:0] put_Data_0_1361;
  reg [8-1:0] put_Key_1_1362;
  reg [1-1:0] put_KeyCompares_1_1363;
  reg [3-1:0] put_KeyCollapse_1_1364;
  reg [8-1:0] put_Data_1_1365;
  reg [8-1:0] put_Key_2_1366;
  reg [1-1:0] put_KeyCompares_2_1367;
  reg [3-1:0] put_KeyCollapse_2_1368;
  reg [8-1:0] put_Data_2_1369;
  reg [8-1:0] put_Key_3_1370;
  reg [1-1:0] put_KeyCompares_3_1371;
  reg [3-1:0] put_KeyCollapse_3_1372;
  reg [8-1:0] put_Data_3_1373;
  reg [1-1:0] put_Found_1374;
  reg [8-1:0] put_Key_1375;
  reg [8-1:0] put_FoundKey_1376;
  reg [8-1:0] put_Data_1377;
  reg [6-1:0] put_BtreeIndex_1378;
  reg [3-1:0] put_StuckIndex_1379;
  reg [1-1:0] put_MergeSuccess_1380;
  reg [6-1:0] put_index_1381;
  reg [3-1:0] put_size_1382;
  reg [1-1:0] put_isLeaf_1383;
  reg [6-1:0] put_nextFree_1384;
  reg [8-1:0] put_Key_0_1385;
  reg [1-1:0] put_KeyCompares_0_1386;
  reg [3-1:0] put_KeyCollapse_0_1387;
  reg [8-1:0] put_Data_0_1388;
  reg [8-1:0] put_Key_1_1389;
  reg [1-1:0] put_KeyCompares_1_1390;
  reg [3-1:0] put_KeyCollapse_1_1391;
  reg [8-1:0] put_Data_1_1392;
  reg [8-1:0] put_Key_2_1393;
  reg [1-1:0] put_KeyCompares_2_1394;
  reg [3-1:0] put_KeyCollapse_2_1395;
  reg [8-1:0] put_Data_2_1396;
  reg [8-1:0] put_Key_3_1397;
  reg [1-1:0] put_KeyCompares_3_1398;
  reg [3-1:0] put_KeyCollapse_3_1399;
  reg [8-1:0] put_Data_3_1400;
  reg [1-1:0] put_Found_1401;
  reg [8-1:0] put_Key_1402;
  reg [8-1:0] put_FoundKey_1403;
  reg [8-1:0] put_Data_1404;
  reg [6-1:0] put_BtreeIndex_1405;
  reg [3-1:0] put_StuckIndex_1406;
  reg [1-1:0] put_MergeSuccess_1407;
  reg [8-1:0] put_childKey_1408;
  reg [6-1:0] put_childData_1409;
  reg [6-1:0] put_indexLeft_1410;
  reg [6-1:0] put_indexRight_1411;
  reg [8-1:0] put_midKey_1412;
  reg [1-1:0] put_success_1413;
  reg [1-1:0] put_test_1414;
  reg [6-1:0] put_next_1415;
  reg [6-1:0] put_root_1416;
  reg [1-1:0] put_isFree_1417;
  reg [6-1:0] put_index_1418;
  reg [3-1:0] put_size_1419;
  reg [1-1:0] put_isLeaf_1420;
  reg [6-1:0] put_nextFree_1421;
  reg [8-1:0] put_Key_0_1422;
  reg [1-1:0] put_KeyCompares_0_1423;
  reg [3-1:0] put_KeyCollapse_0_1424;
  reg [8-1:0] put_Data_0_1425;
  reg [8-1:0] put_Key_1_1426;
  reg [1-1:0] put_KeyCompares_1_1427;
  reg [3-1:0] put_KeyCollapse_1_1428;
  reg [8-1:0] put_Data_1_1429;
  reg [8-1:0] put_Key_2_1430;
  reg [1-1:0] put_KeyCompares_2_1431;
  reg [3-1:0] put_KeyCollapse_2_1432;
  reg [8-1:0] put_Data_2_1433;
  reg [8-1:0] put_Key_3_1434;
  reg [1-1:0] put_KeyCompares_3_1435;
  reg [3-1:0] put_KeyCollapse_3_1436;
  reg [8-1:0] put_Data_3_1437;
  reg [1-1:0] put_Found_1438;
  reg [8-1:0] put_Key_1439;
  reg [8-1:0] put_FoundKey_1440;
  reg [8-1:0] put_Data_1441;
  reg [6-1:0] put_BtreeIndex_1442;
  reg [3-1:0] put_StuckIndex_1443;
  reg [1-1:0] put_MergeSuccess_1444;
  reg [6-1:0] put_index_1445;
  reg [3-1:0] put_size_1446;
  reg [1-1:0] put_isLeaf_1447;
  reg [6-1:0] put_nextFree_1448;
  reg [8-1:0] put_Key_0_1449;
  reg [1-1:0] put_KeyCompares_0_1450;
  reg [3-1:0] put_KeyCollapse_0_1451;
  reg [8-1:0] put_Data_0_1452;
  reg [8-1:0] put_Key_1_1453;
  reg [1-1:0] put_KeyCompares_1_1454;
  reg [3-1:0] put_KeyCollapse_1_1455;
  reg [8-1:0] put_Data_1_1456;
  reg [8-1:0] put_Key_2_1457;
  reg [1-1:0] put_KeyCompares_2_1458;
  reg [3-1:0] put_KeyCollapse_2_1459;
  reg [8-1:0] put_Data_2_1460;
  reg [8-1:0] put_Key_3_1461;
  reg [1-1:0] put_KeyCompares_3_1462;
  reg [3-1:0] put_KeyCollapse_3_1463;
  reg [8-1:0] put_Data_3_1464;
  reg [1-1:0] put_Found_1465;
  reg [8-1:0] put_Key_1466;
  reg [8-1:0] put_FoundKey_1467;
  reg [8-1:0] put_Data_1468;
  reg [6-1:0] put_BtreeIndex_1469;
  reg [3-1:0] put_StuckIndex_1470;
  reg [1-1:0] put_MergeSuccess_1471;
  reg [8-1:0] put_childKey_1472;
  reg [3-1:0] put_leftChild_1473;
  reg [3-1:0] put_rightChild_1474;
  reg [6-1:0] put_childData_1475;
  reg [6-1:0] put_indexLeft_1476;
  reg [6-1:0] put_indexRight_1477;
  reg [8-1:0] put_midKey_1478;
  reg [1-1:0] put_success_1479;
  reg [1-1:0] put_test_1480;
  reg [6-1:0] put_next_1481;
  reg [6-1:0] put_root_1482;
  reg [1-1:0] put_isFree_1483;
  integer put_pc;
  integer put_stop;
  integer put_returnCode;
  integer put_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      put_pc <= 0;
      put_stop <= 0;
      put_returnCode <= 0;
      put_k_0 <= 0;
      put_d_1 <= 0;
      put_i_2 <= 0;
      put_l_3 <= 0;
      put_index_4 <= 0;
      put_size_5 <= 0;
      put_isLeaf_6 <= 0;
      put_nextFree_7 <= 0;
      put_Key_0_8 <= 0;
      put_KeyCompares_0_9 <= 0;
      put_KeyCollapse_0_10 <= 0;
      put_Data_0_11 <= 0;
      put_Key_1_12 <= 0;
      put_KeyCompares_1_13 <= 0;
      put_KeyCollapse_1_14 <= 0;
      put_Data_1_15 <= 0;
      put_Key_2_16 <= 0;
      put_KeyCompares_2_17 <= 0;
      put_KeyCollapse_2_18 <= 0;
      put_Data_2_19 <= 0;
      put_Key_3_20 <= 0;
      put_KeyCompares_3_21 <= 0;
      put_KeyCollapse_3_22 <= 0;
      put_Data_3_23 <= 0;
      put_stuckKeys_1_index_24 <= 0;
      put_stuckKeys_2_index_25 <= 0;
      put_stuckKeys_2_value_26 <= 0;
      put_stuckKeys_2_value_27 <= 0;
      put_stuckKeys_2_value_28 <= 0;
      put_stuckKeys_2_value_29 <= 0;
      put_stuckData_3_index_30 <= 0;
      put_stuckData_4_index_31 <= 0;
      put_stuckData_4_value_32 <= 0;
      put_stuckData_4_value_33 <= 0;
      put_stuckData_4_value_34 <= 0;
      put_stuckData_4_value_35 <= 0;
      put_stuckSize_5_index_36 <= 0;
      put_stuckSize_6_index_37 <= 0;
      put_stuckSize_6_value_38 <= 0;
      put_stuckIsLeaf_7_index_39 <= 0;
      put_stuckIsLeaf_8_index_40 <= 0;
      put_stuckIsLeaf_8_value_41 <= 0;
      put_Found_42 <= 0;
      put_Key_43 <= 0;
      put_FoundKey_44 <= 0;
      put_Data_45 <= 0;
      put_BtreeIndex_46 <= 0;
      put_StuckIndex_47 <= 0;
      put_MergeSuccess_48 <= 0;
      put_index_49 <= 0;
      put_size_50 <= 0;
      put_isLeaf_51 <= 0;
      put_nextFree_52 <= 0;
      put_Key_0_53 <= 0;
      put_KeyCompares_0_54 <= 0;
      put_KeyCollapse_0_55 <= 0;
      put_Data_0_56 <= 0;
      put_Key_1_57 <= 0;
      put_KeyCompares_1_58 <= 0;
      put_KeyCollapse_1_59 <= 0;
      put_Data_1_60 <= 0;
      put_Key_2_61 <= 0;
      put_KeyCompares_2_62 <= 0;
      put_KeyCollapse_2_63 <= 0;
      put_Data_2_64 <= 0;
      put_Key_3_65 <= 0;
      put_KeyCompares_3_66 <= 0;
      put_KeyCollapse_3_67 <= 0;
      put_Data_3_68 <= 0;
      put_Found_69 <= 0;
      put_Key_70 <= 0;
      put_FoundKey_71 <= 0;
      put_Data_72 <= 0;
      put_BtreeIndex_73 <= 0;
      put_StuckIndex_74 <= 0;
      put_MergeSuccess_75 <= 0;
      put_index_76 <= 0;
      put_size_77 <= 0;
      put_isLeaf_78 <= 0;
      put_nextFree_79 <= 0;
      put_Key_0_80 <= 0;
      put_KeyCompares_0_81 <= 0;
      put_KeyCollapse_0_82 <= 0;
      put_Data_0_83 <= 0;
      put_Key_1_84 <= 0;
      put_KeyCompares_1_85 <= 0;
      put_KeyCollapse_1_86 <= 0;
      put_Data_1_87 <= 0;
      put_Key_2_88 <= 0;
      put_KeyCompares_2_89 <= 0;
      put_KeyCollapse_2_90 <= 0;
      put_Data_2_91 <= 0;
      put_Key_3_92 <= 0;
      put_KeyCompares_3_93 <= 0;
      put_KeyCollapse_3_94 <= 0;
      put_Data_3_95 <= 0;
      put_Found_96 <= 0;
      put_Key_97 <= 0;
      put_FoundKey_98 <= 0;
      put_Data_99 <= 0;
      put_BtreeIndex_100 <= 0;
      put_StuckIndex_101 <= 0;
      put_MergeSuccess_102 <= 0;
      put_child_103 <= 0;
      put_parent_104 <= 0;
      put_childInparent_105 <= 0;
      put_found_106 <= 0;
      put_full_107 <= 0;
      put_i_108 <= 0;
      put_notFull_109 <= 0;
      put_index_110 <= 0;
      put_size_111 <= 0;
      put_isLeaf_112 <= 0;
      put_nextFree_113 <= 0;
      put_Key_0_114 <= 0;
      put_KeyCompares_0_115 <= 0;
      put_KeyCollapse_0_116 <= 0;
      put_Data_0_117 <= 0;
      put_Key_1_118 <= 0;
      put_KeyCompares_1_119 <= 0;
      put_KeyCollapse_1_120 <= 0;
      put_Data_1_121 <= 0;
      put_Key_2_122 <= 0;
      put_KeyCompares_2_123 <= 0;
      put_KeyCollapse_2_124 <= 0;
      put_Data_2_125 <= 0;
      put_Key_3_126 <= 0;
      put_KeyCompares_3_127 <= 0;
      put_KeyCollapse_3_128 <= 0;
      put_Data_3_129 <= 0;
      put_Found_130 <= 0;
      put_Key_131 <= 0;
      put_FoundKey_132 <= 0;
      put_Data_133 <= 0;
      put_BtreeIndex_134 <= 0;
      put_StuckIndex_135 <= 0;
      put_MergeSuccess_136 <= 0;
      put_index_137 <= 0;
      put_size_138 <= 0;
      put_isLeaf_139 <= 0;
      put_nextFree_140 <= 0;
      put_Key_0_141 <= 0;
      put_KeyCompares_0_142 <= 0;
      put_KeyCollapse_0_143 <= 0;
      put_Data_0_144 <= 0;
      put_Key_1_145 <= 0;
      put_KeyCompares_1_146 <= 0;
      put_KeyCollapse_1_147 <= 0;
      put_Data_1_148 <= 0;
      put_Key_2_149 <= 0;
      put_KeyCompares_2_150 <= 0;
      put_KeyCollapse_2_151 <= 0;
      put_Data_2_152 <= 0;
      put_Key_3_153 <= 0;
      put_KeyCompares_3_154 <= 0;
      put_KeyCollapse_3_155 <= 0;
      put_Data_3_156 <= 0;
      put_Found_157 <= 0;
      put_Key_158 <= 0;
      put_FoundKey_159 <= 0;
      put_Data_160 <= 0;
      put_BtreeIndex_161 <= 0;
      put_StuckIndex_162 <= 0;
      put_MergeSuccess_163 <= 0;
      put_index_164 <= 0;
      put_size_165 <= 0;
      put_isLeaf_166 <= 0;
      put_nextFree_167 <= 0;
      put_Key_0_168 <= 0;
      put_KeyCompares_0_169 <= 0;
      put_KeyCollapse_0_170 <= 0;
      put_Data_0_171 <= 0;
      put_Key_1_172 <= 0;
      put_KeyCompares_1_173 <= 0;
      put_KeyCollapse_1_174 <= 0;
      put_Data_1_175 <= 0;
      put_Key_2_176 <= 0;
      put_KeyCompares_2_177 <= 0;
      put_KeyCollapse_2_178 <= 0;
      put_Data_2_179 <= 0;
      put_Key_3_180 <= 0;
      put_KeyCompares_3_181 <= 0;
      put_KeyCollapse_3_182 <= 0;
      put_Data_3_183 <= 0;
      put_Found_184 <= 0;
      put_Key_185 <= 0;
      put_FoundKey_186 <= 0;
      put_Data_187 <= 0;
      put_BtreeIndex_188 <= 0;
      put_StuckIndex_189 <= 0;
      put_MergeSuccess_190 <= 0;
      put_indexLeft_191 <= 0;
      put_indexRight_192 <= 0;
      put_midKey_193 <= 0;
      put_freeNext_9_index_194 <= 0;
      put_freeNext_10_index_195 <= 0;
      put_freeNext_10_value_196 <= 0;
      put_stuckIsFree_11_index_197 <= 0;
      put_stuckIsFree_11_value_198 <= 0;
      put_root_199 <= 0;
      put_next_200 <= 0;
      put_isLeaf_201 <= 0;
      put_isFree_202 <= 0;
      put_root_203 <= 0;
      put_next_204 <= 0;
      put_isLeaf_205 <= 0;
      put_isFree_206 <= 0;
      put_i_207 <= 0;
      put_notFull_208 <= 0;
      put_index_209 <= 0;
      put_size_210 <= 0;
      put_isLeaf_211 <= 0;
      put_nextFree_212 <= 0;
      put_Key_0_213 <= 0;
      put_KeyCompares_0_214 <= 0;
      put_KeyCollapse_0_215 <= 0;
      put_Data_0_216 <= 0;
      put_Key_1_217 <= 0;
      put_KeyCompares_1_218 <= 0;
      put_KeyCollapse_1_219 <= 0;
      put_Data_1_220 <= 0;
      put_Key_2_221 <= 0;
      put_KeyCompares_2_222 <= 0;
      put_KeyCollapse_2_223 <= 0;
      put_Data_2_224 <= 0;
      put_Key_3_225 <= 0;
      put_KeyCompares_3_226 <= 0;
      put_KeyCollapse_3_227 <= 0;
      put_Data_3_228 <= 0;
      put_Found_229 <= 0;
      put_Key_230 <= 0;
      put_FoundKey_231 <= 0;
      put_Data_232 <= 0;
      put_BtreeIndex_233 <= 0;
      put_StuckIndex_234 <= 0;
      put_MergeSuccess_235 <= 0;
      put_index_236 <= 0;
      put_size_237 <= 0;
      put_isLeaf_238 <= 0;
      put_nextFree_239 <= 0;
      put_Key_0_240 <= 0;
      put_KeyCompares_0_241 <= 0;
      put_KeyCollapse_0_242 <= 0;
      put_Data_0_243 <= 0;
      put_Key_1_244 <= 0;
      put_KeyCompares_1_245 <= 0;
      put_KeyCollapse_1_246 <= 0;
      put_Data_1_247 <= 0;
      put_Key_2_248 <= 0;
      put_KeyCompares_2_249 <= 0;
      put_KeyCollapse_2_250 <= 0;
      put_Data_2_251 <= 0;
      put_Key_3_252 <= 0;
      put_KeyCompares_3_253 <= 0;
      put_KeyCollapse_3_254 <= 0;
      put_Data_3_255 <= 0;
      put_Found_256 <= 0;
      put_Key_257 <= 0;
      put_FoundKey_258 <= 0;
      put_Data_259 <= 0;
      put_BtreeIndex_260 <= 0;
      put_StuckIndex_261 <= 0;
      put_MergeSuccess_262 <= 0;
      put_index_263 <= 0;
      put_size_264 <= 0;
      put_isLeaf_265 <= 0;
      put_nextFree_266 <= 0;
      put_Key_0_267 <= 0;
      put_KeyCompares_0_268 <= 0;
      put_KeyCollapse_0_269 <= 0;
      put_Data_0_270 <= 0;
      put_Key_1_271 <= 0;
      put_KeyCompares_1_272 <= 0;
      put_KeyCollapse_1_273 <= 0;
      put_Data_1_274 <= 0;
      put_Key_2_275 <= 0;
      put_KeyCompares_2_276 <= 0;
      put_KeyCollapse_2_277 <= 0;
      put_Data_2_278 <= 0;
      put_Key_3_279 <= 0;
      put_KeyCompares_3_280 <= 0;
      put_KeyCollapse_3_281 <= 0;
      put_Data_3_282 <= 0;
      put_Found_283 <= 0;
      put_Key_284 <= 0;
      put_FoundKey_285 <= 0;
      put_Data_286 <= 0;
      put_BtreeIndex_287 <= 0;
      put_StuckIndex_288 <= 0;
      put_MergeSuccess_289 <= 0;
      put_indexLeft_290 <= 0;
      put_indexRight_291 <= 0;
      put_midKey_292 <= 0;
      put_root_293 <= 0;
      put_next_294 <= 0;
      put_isLeaf_295 <= 0;
      put_isFree_296 <= 0;
      put_root_297 <= 0;
      put_next_298 <= 0;
      put_isLeaf_299 <= 0;
      put_isFree_300 <= 0;
      put_index_301 <= 0;
      put_size_302 <= 0;
      put_isLeaf_303 <= 0;
      put_nextFree_304 <= 0;
      put_Key_0_305 <= 0;
      put_KeyCompares_0_306 <= 0;
      put_KeyCollapse_0_307 <= 0;
      put_Data_0_308 <= 0;
      put_Key_1_309 <= 0;
      put_KeyCompares_1_310 <= 0;
      put_KeyCollapse_1_311 <= 0;
      put_Data_1_312 <= 0;
      put_Key_2_313 <= 0;
      put_KeyCompares_2_314 <= 0;
      put_KeyCollapse_2_315 <= 0;
      put_Data_2_316 <= 0;
      put_Key_3_317 <= 0;
      put_KeyCompares_3_318 <= 0;
      put_KeyCollapse_3_319 <= 0;
      put_Data_3_320 <= 0;
      put_Found_321 <= 0;
      put_Key_322 <= 0;
      put_FoundKey_323 <= 0;
      put_Data_324 <= 0;
      put_BtreeIndex_325 <= 0;
      put_StuckIndex_326 <= 0;
      put_MergeSuccess_327 <= 0;
      put_index_328 <= 0;
      put_size_329 <= 0;
      put_isLeaf_330 <= 0;
      put_nextFree_331 <= 0;
      put_Key_0_332 <= 0;
      put_KeyCompares_0_333 <= 0;
      put_KeyCollapse_0_334 <= 0;
      put_Data_0_335 <= 0;
      put_Key_1_336 <= 0;
      put_KeyCompares_1_337 <= 0;
      put_KeyCollapse_1_338 <= 0;
      put_Data_1_339 <= 0;
      put_Key_2_340 <= 0;
      put_KeyCompares_2_341 <= 0;
      put_KeyCollapse_2_342 <= 0;
      put_Data_2_343 <= 0;
      put_Key_3_344 <= 0;
      put_KeyCompares_3_345 <= 0;
      put_KeyCollapse_3_346 <= 0;
      put_Data_3_347 <= 0;
      put_Found_348 <= 0;
      put_Key_349 <= 0;
      put_FoundKey_350 <= 0;
      put_Data_351 <= 0;
      put_BtreeIndex_352 <= 0;
      put_StuckIndex_353 <= 0;
      put_MergeSuccess_354 <= 0;
      put_index_355 <= 0;
      put_size_356 <= 0;
      put_isLeaf_357 <= 0;
      put_nextFree_358 <= 0;
      put_Key_0_359 <= 0;
      put_KeyCompares_0_360 <= 0;
      put_KeyCollapse_0_361 <= 0;
      put_Data_0_362 <= 0;
      put_Key_1_363 <= 0;
      put_KeyCompares_1_364 <= 0;
      put_KeyCollapse_1_365 <= 0;
      put_Data_1_366 <= 0;
      put_Key_2_367 <= 0;
      put_KeyCompares_2_368 <= 0;
      put_KeyCollapse_2_369 <= 0;
      put_Data_2_370 <= 0;
      put_Key_3_371 <= 0;
      put_KeyCompares_3_372 <= 0;
      put_KeyCollapse_3_373 <= 0;
      put_Data_3_374 <= 0;
      put_Found_375 <= 0;
      put_Key_376 <= 0;
      put_FoundKey_377 <= 0;
      put_Data_378 <= 0;
      put_BtreeIndex_379 <= 0;
      put_StuckIndex_380 <= 0;
      put_MergeSuccess_381 <= 0;
      put_index_382 <= 0;
      put_size_383 <= 0;
      put_isLeaf_384 <= 0;
      put_nextFree_385 <= 0;
      put_Key_0_386 <= 0;
      put_KeyCompares_0_387 <= 0;
      put_KeyCollapse_0_388 <= 0;
      put_Data_0_389 <= 0;
      put_Key_1_390 <= 0;
      put_KeyCompares_1_391 <= 0;
      put_KeyCollapse_1_392 <= 0;
      put_Data_1_393 <= 0;
      put_Key_2_394 <= 0;
      put_KeyCompares_2_395 <= 0;
      put_KeyCollapse_2_396 <= 0;
      put_Data_2_397 <= 0;
      put_Key_3_398 <= 0;
      put_KeyCompares_3_399 <= 0;
      put_KeyCollapse_3_400 <= 0;
      put_Data_3_401 <= 0;
      put_Found_402 <= 0;
      put_Key_403 <= 0;
      put_FoundKey_404 <= 0;
      put_Data_405 <= 0;
      put_BtreeIndex_406 <= 0;
      put_StuckIndex_407 <= 0;
      put_MergeSuccess_408 <= 0;
      put_childKey_409 <= 0;
      put_childData_410 <= 0;
      put_indexLeft_411 <= 0;
      put_indexRight_412 <= 0;
      put_midKey_413 <= 0;
      put_root_414 <= 0;
      put_next_415 <= 0;
      put_isLeaf_416 <= 0;
      put_isFree_417 <= 0;
      put_index_418 <= 0;
      put_size_419 <= 0;
      put_isLeaf_420 <= 0;
      put_nextFree_421 <= 0;
      put_Key_0_422 <= 0;
      put_KeyCompares_0_423 <= 0;
      put_KeyCollapse_0_424 <= 0;
      put_Data_0_425 <= 0;
      put_Key_1_426 <= 0;
      put_KeyCompares_1_427 <= 0;
      put_KeyCollapse_1_428 <= 0;
      put_Data_1_429 <= 0;
      put_Key_2_430 <= 0;
      put_KeyCompares_2_431 <= 0;
      put_KeyCollapse_2_432 <= 0;
      put_Data_2_433 <= 0;
      put_Key_3_434 <= 0;
      put_KeyCompares_3_435 <= 0;
      put_KeyCollapse_3_436 <= 0;
      put_Data_3_437 <= 0;
      put_Found_438 <= 0;
      put_Key_439 <= 0;
      put_FoundKey_440 <= 0;
      put_Data_441 <= 0;
      put_BtreeIndex_442 <= 0;
      put_StuckIndex_443 <= 0;
      put_MergeSuccess_444 <= 0;
      put_index_445 <= 0;
      put_size_446 <= 0;
      put_isLeaf_447 <= 0;
      put_nextFree_448 <= 0;
      put_Key_0_449 <= 0;
      put_KeyCompares_0_450 <= 0;
      put_KeyCollapse_0_451 <= 0;
      put_Data_0_452 <= 0;
      put_Key_1_453 <= 0;
      put_KeyCompares_1_454 <= 0;
      put_KeyCollapse_1_455 <= 0;
      put_Data_1_456 <= 0;
      put_Key_2_457 <= 0;
      put_KeyCompares_2_458 <= 0;
      put_KeyCollapse_2_459 <= 0;
      put_Data_2_460 <= 0;
      put_Key_3_461 <= 0;
      put_KeyCompares_3_462 <= 0;
      put_KeyCollapse_3_463 <= 0;
      put_Data_3_464 <= 0;
      put_Found_465 <= 0;
      put_Key_466 <= 0;
      put_FoundKey_467 <= 0;
      put_Data_468 <= 0;
      put_BtreeIndex_469 <= 0;
      put_StuckIndex_470 <= 0;
      put_MergeSuccess_471 <= 0;
      put_index_472 <= 0;
      put_size_473 <= 0;
      put_isLeaf_474 <= 0;
      put_nextFree_475 <= 0;
      put_Key_0_476 <= 0;
      put_KeyCompares_0_477 <= 0;
      put_KeyCollapse_0_478 <= 0;
      put_Data_0_479 <= 0;
      put_Key_1_480 <= 0;
      put_KeyCompares_1_481 <= 0;
      put_KeyCollapse_1_482 <= 0;
      put_Data_1_483 <= 0;
      put_Key_2_484 <= 0;
      put_KeyCompares_2_485 <= 0;
      put_KeyCollapse_2_486 <= 0;
      put_Data_2_487 <= 0;
      put_Key_3_488 <= 0;
      put_KeyCompares_3_489 <= 0;
      put_KeyCollapse_3_490 <= 0;
      put_Data_3_491 <= 0;
      put_Found_492 <= 0;
      put_Key_493 <= 0;
      put_FoundKey_494 <= 0;
      put_Data_495 <= 0;
      put_BtreeIndex_496 <= 0;
      put_StuckIndex_497 <= 0;
      put_MergeSuccess_498 <= 0;
      put_childIndex_499 <= 0;
      put_leftIndex_500 <= 0;
      put_midKey_501 <= 0;
      put_root_502 <= 0;
      put_next_503 <= 0;
      put_isLeaf_504 <= 0;
      put_isFree_505 <= 0;
      put_i_506 <= 0;
      put_notFull_507 <= 0;
      put_index_508 <= 0;
      put_size_509 <= 0;
      put_isLeaf_510 <= 0;
      put_nextFree_511 <= 0;
      put_Key_0_512 <= 0;
      put_KeyCompares_0_513 <= 0;
      put_KeyCollapse_0_514 <= 0;
      put_Data_0_515 <= 0;
      put_Key_1_516 <= 0;
      put_KeyCompares_1_517 <= 0;
      put_KeyCollapse_1_518 <= 0;
      put_Data_1_519 <= 0;
      put_Key_2_520 <= 0;
      put_KeyCompares_2_521 <= 0;
      put_KeyCollapse_2_522 <= 0;
      put_Data_2_523 <= 0;
      put_Key_3_524 <= 0;
      put_KeyCompares_3_525 <= 0;
      put_KeyCollapse_3_526 <= 0;
      put_Data_3_527 <= 0;
      put_Found_528 <= 0;
      put_Key_529 <= 0;
      put_FoundKey_530 <= 0;
      put_Data_531 <= 0;
      put_BtreeIndex_532 <= 0;
      put_StuckIndex_533 <= 0;
      put_MergeSuccess_534 <= 0;
      put_index_535 <= 0;
      put_size_536 <= 0;
      put_isLeaf_537 <= 0;
      put_nextFree_538 <= 0;
      put_Key_0_539 <= 0;
      put_KeyCompares_0_540 <= 0;
      put_KeyCollapse_0_541 <= 0;
      put_Data_0_542 <= 0;
      put_Key_1_543 <= 0;
      put_KeyCompares_1_544 <= 0;
      put_KeyCollapse_1_545 <= 0;
      put_Data_1_546 <= 0;
      put_Key_2_547 <= 0;
      put_KeyCompares_2_548 <= 0;
      put_KeyCollapse_2_549 <= 0;
      put_Data_2_550 <= 0;
      put_Key_3_551 <= 0;
      put_KeyCompares_3_552 <= 0;
      put_KeyCollapse_3_553 <= 0;
      put_Data_3_554 <= 0;
      put_Found_555 <= 0;
      put_Key_556 <= 0;
      put_FoundKey_557 <= 0;
      put_Data_558 <= 0;
      put_BtreeIndex_559 <= 0;
      put_StuckIndex_560 <= 0;
      put_MergeSuccess_561 <= 0;
      put_index_562 <= 0;
      put_size_563 <= 0;
      put_isLeaf_564 <= 0;
      put_nextFree_565 <= 0;
      put_Key_0_566 <= 0;
      put_KeyCompares_0_567 <= 0;
      put_KeyCollapse_0_568 <= 0;
      put_Data_0_569 <= 0;
      put_Key_1_570 <= 0;
      put_KeyCompares_1_571 <= 0;
      put_KeyCollapse_1_572 <= 0;
      put_Data_1_573 <= 0;
      put_Key_2_574 <= 0;
      put_KeyCompares_2_575 <= 0;
      put_KeyCollapse_2_576 <= 0;
      put_Data_2_577 <= 0;
      put_Key_3_578 <= 0;
      put_KeyCompares_3_579 <= 0;
      put_KeyCollapse_3_580 <= 0;
      put_Data_3_581 <= 0;
      put_Found_582 <= 0;
      put_Key_583 <= 0;
      put_FoundKey_584 <= 0;
      put_Data_585 <= 0;
      put_BtreeIndex_586 <= 0;
      put_StuckIndex_587 <= 0;
      put_MergeSuccess_588 <= 0;
      put_index_589 <= 0;
      put_size_590 <= 0;
      put_isLeaf_591 <= 0;
      put_nextFree_592 <= 0;
      put_Key_0_593 <= 0;
      put_KeyCompares_0_594 <= 0;
      put_KeyCollapse_0_595 <= 0;
      put_Data_0_596 <= 0;
      put_Key_1_597 <= 0;
      put_KeyCompares_1_598 <= 0;
      put_KeyCollapse_1_599 <= 0;
      put_Data_1_600 <= 0;
      put_Key_2_601 <= 0;
      put_KeyCompares_2_602 <= 0;
      put_KeyCollapse_2_603 <= 0;
      put_Data_2_604 <= 0;
      put_Key_3_605 <= 0;
      put_KeyCompares_3_606 <= 0;
      put_KeyCollapse_3_607 <= 0;
      put_Data_3_608 <= 0;
      put_Found_609 <= 0;
      put_Key_610 <= 0;
      put_FoundKey_611 <= 0;
      put_Data_612 <= 0;
      put_BtreeIndex_613 <= 0;
      put_StuckIndex_614 <= 0;
      put_MergeSuccess_615 <= 0;
      put_childKey_616 <= 0;
      put_childData_617 <= 0;
      put_indexLeft_618 <= 0;
      put_indexRight_619 <= 0;
      put_midKey_620 <= 0;
      put_root_621 <= 0;
      put_next_622 <= 0;
      put_isLeaf_623 <= 0;
      put_isFree_624 <= 0;
      put_index_625 <= 0;
      put_size_626 <= 0;
      put_isLeaf_627 <= 0;
      put_nextFree_628 <= 0;
      put_Key_0_629 <= 0;
      put_KeyCompares_0_630 <= 0;
      put_KeyCollapse_0_631 <= 0;
      put_Data_0_632 <= 0;
      put_Key_1_633 <= 0;
      put_KeyCompares_1_634 <= 0;
      put_KeyCollapse_1_635 <= 0;
      put_Data_1_636 <= 0;
      put_Key_2_637 <= 0;
      put_KeyCompares_2_638 <= 0;
      put_KeyCollapse_2_639 <= 0;
      put_Data_2_640 <= 0;
      put_Key_3_641 <= 0;
      put_KeyCompares_3_642 <= 0;
      put_KeyCollapse_3_643 <= 0;
      put_Data_3_644 <= 0;
      put_Found_645 <= 0;
      put_Key_646 <= 0;
      put_FoundKey_647 <= 0;
      put_Data_648 <= 0;
      put_BtreeIndex_649 <= 0;
      put_StuckIndex_650 <= 0;
      put_MergeSuccess_651 <= 0;
      put_index_652 <= 0;
      put_size_653 <= 0;
      put_isLeaf_654 <= 0;
      put_nextFree_655 <= 0;
      put_Key_0_656 <= 0;
      put_KeyCompares_0_657 <= 0;
      put_KeyCollapse_0_658 <= 0;
      put_Data_0_659 <= 0;
      put_Key_1_660 <= 0;
      put_KeyCompares_1_661 <= 0;
      put_KeyCollapse_1_662 <= 0;
      put_Data_1_663 <= 0;
      put_Key_2_664 <= 0;
      put_KeyCompares_2_665 <= 0;
      put_KeyCollapse_2_666 <= 0;
      put_Data_2_667 <= 0;
      put_Key_3_668 <= 0;
      put_KeyCompares_3_669 <= 0;
      put_KeyCollapse_3_670 <= 0;
      put_Data_3_671 <= 0;
      put_Found_672 <= 0;
      put_Key_673 <= 0;
      put_FoundKey_674 <= 0;
      put_Data_675 <= 0;
      put_BtreeIndex_676 <= 0;
      put_StuckIndex_677 <= 0;
      put_MergeSuccess_678 <= 0;
      put_index_679 <= 0;
      put_size_680 <= 0;
      put_isLeaf_681 <= 0;
      put_nextFree_682 <= 0;
      put_Key_0_683 <= 0;
      put_KeyCompares_0_684 <= 0;
      put_KeyCollapse_0_685 <= 0;
      put_Data_0_686 <= 0;
      put_Key_1_687 <= 0;
      put_KeyCompares_1_688 <= 0;
      put_KeyCollapse_1_689 <= 0;
      put_Data_1_690 <= 0;
      put_Key_2_691 <= 0;
      put_KeyCompares_2_692 <= 0;
      put_KeyCollapse_2_693 <= 0;
      put_Data_2_694 <= 0;
      put_Key_3_695 <= 0;
      put_KeyCompares_3_696 <= 0;
      put_KeyCollapse_3_697 <= 0;
      put_Data_3_698 <= 0;
      put_Found_699 <= 0;
      put_Key_700 <= 0;
      put_FoundKey_701 <= 0;
      put_Data_702 <= 0;
      put_BtreeIndex_703 <= 0;
      put_StuckIndex_704 <= 0;
      put_MergeSuccess_705 <= 0;
      put_index_706 <= 0;
      put_size_707 <= 0;
      put_isLeaf_708 <= 0;
      put_nextFree_709 <= 0;
      put_Key_0_710 <= 0;
      put_KeyCompares_0_711 <= 0;
      put_KeyCollapse_0_712 <= 0;
      put_Data_0_713 <= 0;
      put_Key_1_714 <= 0;
      put_KeyCompares_1_715 <= 0;
      put_KeyCollapse_1_716 <= 0;
      put_Data_1_717 <= 0;
      put_Key_2_718 <= 0;
      put_KeyCompares_2_719 <= 0;
      put_KeyCollapse_2_720 <= 0;
      put_Data_2_721 <= 0;
      put_Key_3_722 <= 0;
      put_KeyCompares_3_723 <= 0;
      put_KeyCollapse_3_724 <= 0;
      put_Data_3_725 <= 0;
      put_Found_726 <= 0;
      put_Key_727 <= 0;
      put_FoundKey_728 <= 0;
      put_Data_729 <= 0;
      put_BtreeIndex_730 <= 0;
      put_StuckIndex_731 <= 0;
      put_MergeSuccess_732 <= 0;
      put_childKey_733 <= 0;
      put_childData_734 <= 0;
      put_indexLeft_735 <= 0;
      put_indexRight_736 <= 0;
      put_midKey_737 <= 0;
      put_root_738 <= 0;
      put_next_739 <= 0;
      put_isLeaf_740 <= 0;
      put_isFree_741 <= 0;
      put_index_742 <= 0;
      put_size_743 <= 0;
      put_isLeaf_744 <= 0;
      put_nextFree_745 <= 0;
      put_Key_0_746 <= 0;
      put_KeyCompares_0_747 <= 0;
      put_KeyCollapse_0_748 <= 0;
      put_Data_0_749 <= 0;
      put_Key_1_750 <= 0;
      put_KeyCompares_1_751 <= 0;
      put_KeyCollapse_1_752 <= 0;
      put_Data_1_753 <= 0;
      put_Key_2_754 <= 0;
      put_KeyCompares_2_755 <= 0;
      put_KeyCollapse_2_756 <= 0;
      put_Data_2_757 <= 0;
      put_Key_3_758 <= 0;
      put_KeyCompares_3_759 <= 0;
      put_KeyCollapse_3_760 <= 0;
      put_Data_3_761 <= 0;
      put_Found_762 <= 0;
      put_Key_763 <= 0;
      put_FoundKey_764 <= 0;
      put_Data_765 <= 0;
      put_BtreeIndex_766 <= 0;
      put_StuckIndex_767 <= 0;
      put_MergeSuccess_768 <= 0;
      put_position_769 <= 0;
      put_index_770 <= 0;
      put_index1_771 <= 0;
      put_within_772 <= 0;
      put_isLeaf_773 <= 0;
      put_index_774 <= 0;
      put_size_775 <= 0;
      put_isLeaf_776 <= 0;
      put_nextFree_777 <= 0;
      put_Key_0_778 <= 0;
      put_KeyCompares_0_779 <= 0;
      put_KeyCollapse_0_780 <= 0;
      put_Data_0_781 <= 0;
      put_Key_1_782 <= 0;
      put_KeyCompares_1_783 <= 0;
      put_KeyCollapse_1_784 <= 0;
      put_Data_1_785 <= 0;
      put_Key_2_786 <= 0;
      put_KeyCompares_2_787 <= 0;
      put_KeyCollapse_2_788 <= 0;
      put_Data_2_789 <= 0;
      put_Key_3_790 <= 0;
      put_KeyCompares_3_791 <= 0;
      put_KeyCollapse_3_792 <= 0;
      put_Data_3_793 <= 0;
      put_Found_794 <= 0;
      put_Key_795 <= 0;
      put_FoundKey_796 <= 0;
      put_Data_797 <= 0;
      put_BtreeIndex_798 <= 0;
      put_StuckIndex_799 <= 0;
      put_MergeSuccess_800 <= 0;
      put_index_801 <= 0;
      put_size_802 <= 0;
      put_isLeaf_803 <= 0;
      put_nextFree_804 <= 0;
      put_Key_0_805 <= 0;
      put_KeyCompares_0_806 <= 0;
      put_KeyCollapse_0_807 <= 0;
      put_Data_0_808 <= 0;
      put_Key_1_809 <= 0;
      put_KeyCompares_1_810 <= 0;
      put_KeyCollapse_1_811 <= 0;
      put_Data_1_812 <= 0;
      put_Key_2_813 <= 0;
      put_KeyCompares_2_814 <= 0;
      put_KeyCollapse_2_815 <= 0;
      put_Data_2_816 <= 0;
      put_Key_3_817 <= 0;
      put_KeyCompares_3_818 <= 0;
      put_KeyCollapse_3_819 <= 0;
      put_Data_3_820 <= 0;
      put_Found_821 <= 0;
      put_Key_822 <= 0;
      put_FoundKey_823 <= 0;
      put_Data_824 <= 0;
      put_BtreeIndex_825 <= 0;
      put_StuckIndex_826 <= 0;
      put_MergeSuccess_827 <= 0;
      put_index_828 <= 0;
      put_size_829 <= 0;
      put_isLeaf_830 <= 0;
      put_nextFree_831 <= 0;
      put_Key_0_832 <= 0;
      put_KeyCompares_0_833 <= 0;
      put_KeyCollapse_0_834 <= 0;
      put_Data_0_835 <= 0;
      put_Key_1_836 <= 0;
      put_KeyCompares_1_837 <= 0;
      put_KeyCollapse_1_838 <= 0;
      put_Data_1_839 <= 0;
      put_Key_2_840 <= 0;
      put_KeyCompares_2_841 <= 0;
      put_KeyCollapse_2_842 <= 0;
      put_Data_2_843 <= 0;
      put_Key_3_844 <= 0;
      put_KeyCompares_3_845 <= 0;
      put_KeyCollapse_3_846 <= 0;
      put_Data_3_847 <= 0;
      put_Found_848 <= 0;
      put_Key_849 <= 0;
      put_FoundKey_850 <= 0;
      put_Data_851 <= 0;
      put_BtreeIndex_852 <= 0;
      put_StuckIndex_853 <= 0;
      put_MergeSuccess_854 <= 0;
      put_childKey_855 <= 0;
      put_childData_856 <= 0;
      put_indexLeft_857 <= 0;
      put_indexRight_858 <= 0;
      put_midKey_859 <= 0;
      put_success_860 <= 0;
      put_test_861 <= 0;
      put_next_862 <= 0;
      put_root_863 <= 0;
      put_isFree_864 <= 0;
      put_next_865 <= 0;
      put_root_866 <= 0;
      put_isFree_867 <= 0;
      put_index_868 <= 0;
      put_size_869 <= 0;
      put_isLeaf_870 <= 0;
      put_nextFree_871 <= 0;
      put_Key_0_872 <= 0;
      put_KeyCompares_0_873 <= 0;
      put_KeyCollapse_0_874 <= 0;
      put_Data_0_875 <= 0;
      put_Key_1_876 <= 0;
      put_KeyCompares_1_877 <= 0;
      put_KeyCollapse_1_878 <= 0;
      put_Data_1_879 <= 0;
      put_Key_2_880 <= 0;
      put_KeyCompares_2_881 <= 0;
      put_KeyCollapse_2_882 <= 0;
      put_Data_2_883 <= 0;
      put_Key_3_884 <= 0;
      put_KeyCompares_3_885 <= 0;
      put_KeyCollapse_3_886 <= 0;
      put_Data_3_887 <= 0;
      put_Found_888 <= 0;
      put_Key_889 <= 0;
      put_FoundKey_890 <= 0;
      put_Data_891 <= 0;
      put_BtreeIndex_892 <= 0;
      put_StuckIndex_893 <= 0;
      put_MergeSuccess_894 <= 0;
      put_index_895 <= 0;
      put_size_896 <= 0;
      put_isLeaf_897 <= 0;
      put_nextFree_898 <= 0;
      put_Key_0_899 <= 0;
      put_KeyCompares_0_900 <= 0;
      put_KeyCollapse_0_901 <= 0;
      put_Data_0_902 <= 0;
      put_Key_1_903 <= 0;
      put_KeyCompares_1_904 <= 0;
      put_KeyCollapse_1_905 <= 0;
      put_Data_1_906 <= 0;
      put_Key_2_907 <= 0;
      put_KeyCompares_2_908 <= 0;
      put_KeyCollapse_2_909 <= 0;
      put_Data_2_910 <= 0;
      put_Key_3_911 <= 0;
      put_KeyCompares_3_912 <= 0;
      put_KeyCollapse_3_913 <= 0;
      put_Data_3_914 <= 0;
      put_Found_915 <= 0;
      put_Key_916 <= 0;
      put_FoundKey_917 <= 0;
      put_Data_918 <= 0;
      put_BtreeIndex_919 <= 0;
      put_StuckIndex_920 <= 0;
      put_MergeSuccess_921 <= 0;
      put_index_922 <= 0;
      put_size_923 <= 0;
      put_isLeaf_924 <= 0;
      put_nextFree_925 <= 0;
      put_Key_0_926 <= 0;
      put_KeyCompares_0_927 <= 0;
      put_KeyCollapse_0_928 <= 0;
      put_Data_0_929 <= 0;
      put_Key_1_930 <= 0;
      put_KeyCompares_1_931 <= 0;
      put_KeyCollapse_1_932 <= 0;
      put_Data_1_933 <= 0;
      put_Key_2_934 <= 0;
      put_KeyCompares_2_935 <= 0;
      put_KeyCollapse_2_936 <= 0;
      put_Data_2_937 <= 0;
      put_Key_3_938 <= 0;
      put_KeyCompares_3_939 <= 0;
      put_KeyCollapse_3_940 <= 0;
      put_Data_3_941 <= 0;
      put_Found_942 <= 0;
      put_Key_943 <= 0;
      put_FoundKey_944 <= 0;
      put_Data_945 <= 0;
      put_BtreeIndex_946 <= 0;
      put_StuckIndex_947 <= 0;
      put_MergeSuccess_948 <= 0;
      put_childKey_949 <= 0;
      put_leftChild_950 <= 0;
      put_rightChild_951 <= 0;
      put_childData_952 <= 0;
      put_indexLeft_953 <= 0;
      put_indexRight_954 <= 0;
      put_midKey_955 <= 0;
      put_success_956 <= 0;
      put_test_957 <= 0;
      put_next_958 <= 0;
      put_root_959 <= 0;
      put_isFree_960 <= 0;
      put_next_961 <= 0;
      put_root_962 <= 0;
      put_isFree_963 <= 0;
      put_index_964 <= 0;
      put_size_965 <= 0;
      put_isLeaf_966 <= 0;
      put_nextFree_967 <= 0;
      put_Key_0_968 <= 0;
      put_KeyCompares_0_969 <= 0;
      put_KeyCollapse_0_970 <= 0;
      put_Data_0_971 <= 0;
      put_Key_1_972 <= 0;
      put_KeyCompares_1_973 <= 0;
      put_KeyCollapse_1_974 <= 0;
      put_Data_1_975 <= 0;
      put_Key_2_976 <= 0;
      put_KeyCompares_2_977 <= 0;
      put_KeyCollapse_2_978 <= 0;
      put_Data_2_979 <= 0;
      put_Key_3_980 <= 0;
      put_KeyCompares_3_981 <= 0;
      put_KeyCollapse_3_982 <= 0;
      put_Data_3_983 <= 0;
      put_Found_984 <= 0;
      put_Key_985 <= 0;
      put_FoundKey_986 <= 0;
      put_Data_987 <= 0;
      put_BtreeIndex_988 <= 0;
      put_StuckIndex_989 <= 0;
      put_MergeSuccess_990 <= 0;
      put_index_991 <= 0;
      put_size_992 <= 0;
      put_isLeaf_993 <= 0;
      put_nextFree_994 <= 0;
      put_Key_0_995 <= 0;
      put_KeyCompares_0_996 <= 0;
      put_KeyCollapse_0_997 <= 0;
      put_Data_0_998 <= 0;
      put_Key_1_999 <= 0;
      put_KeyCompares_1_1000 <= 0;
      put_KeyCollapse_1_1001 <= 0;
      put_Data_1_1002 <= 0;
      put_Key_2_1003 <= 0;
      put_KeyCompares_2_1004 <= 0;
      put_KeyCollapse_2_1005 <= 0;
      put_Data_2_1006 <= 0;
      put_Key_3_1007 <= 0;
      put_KeyCompares_3_1008 <= 0;
      put_KeyCollapse_3_1009 <= 0;
      put_Data_3_1010 <= 0;
      put_Found_1011 <= 0;
      put_Key_1012 <= 0;
      put_FoundKey_1013 <= 0;
      put_Data_1014 <= 0;
      put_BtreeIndex_1015 <= 0;
      put_StuckIndex_1016 <= 0;
      put_MergeSuccess_1017 <= 0;
      put_childKey_1018 <= 0;
      put_size_1019 <= 0;
      put_childData_1020 <= 0;
      put_indexLeft_1021 <= 0;
      put_indexRight_1022 <= 0;
      put_midKey_1023 <= 0;
      put_success_1024 <= 0;
      put_test_1025 <= 0;
      put_next_1026 <= 0;
      put_root_1027 <= 0;
      put_isFree_1028 <= 0;
      put_index_1029 <= 0;
      put_size_1030 <= 0;
      put_isLeaf_1031 <= 0;
      put_nextFree_1032 <= 0;
      put_Key_0_1033 <= 0;
      put_KeyCompares_0_1034 <= 0;
      put_KeyCollapse_0_1035 <= 0;
      put_Data_0_1036 <= 0;
      put_Key_1_1037 <= 0;
      put_KeyCompares_1_1038 <= 0;
      put_KeyCollapse_1_1039 <= 0;
      put_Data_1_1040 <= 0;
      put_Key_2_1041 <= 0;
      put_KeyCompares_2_1042 <= 0;
      put_KeyCollapse_2_1043 <= 0;
      put_Data_2_1044 <= 0;
      put_Key_3_1045 <= 0;
      put_KeyCompares_3_1046 <= 0;
      put_KeyCollapse_3_1047 <= 0;
      put_Data_3_1048 <= 0;
      put_Found_1049 <= 0;
      put_Key_1050 <= 0;
      put_FoundKey_1051 <= 0;
      put_Data_1052 <= 0;
      put_BtreeIndex_1053 <= 0;
      put_StuckIndex_1054 <= 0;
      put_MergeSuccess_1055 <= 0;
      put_index_1056 <= 0;
      put_size_1057 <= 0;
      put_isLeaf_1058 <= 0;
      put_nextFree_1059 <= 0;
      put_Key_0_1060 <= 0;
      put_KeyCompares_0_1061 <= 0;
      put_KeyCollapse_0_1062 <= 0;
      put_Data_0_1063 <= 0;
      put_Key_1_1064 <= 0;
      put_KeyCompares_1_1065 <= 0;
      put_KeyCollapse_1_1066 <= 0;
      put_Data_1_1067 <= 0;
      put_Key_2_1068 <= 0;
      put_KeyCompares_2_1069 <= 0;
      put_KeyCollapse_2_1070 <= 0;
      put_Data_2_1071 <= 0;
      put_Key_3_1072 <= 0;
      put_KeyCompares_3_1073 <= 0;
      put_KeyCollapse_3_1074 <= 0;
      put_Data_3_1075 <= 0;
      put_Found_1076 <= 0;
      put_Key_1077 <= 0;
      put_FoundKey_1078 <= 0;
      put_Data_1079 <= 0;
      put_BtreeIndex_1080 <= 0;
      put_StuckIndex_1081 <= 0;
      put_MergeSuccess_1082 <= 0;
      put_childKey_1083 <= 0;
      put_size_1084 <= 0;
      put_childData_1085 <= 0;
      put_indexLeft_1086 <= 0;
      put_indexRight_1087 <= 0;
      put_midKey_1088 <= 0;
      put_success_1089 <= 0;
      put_test_1090 <= 0;
      put_next_1091 <= 0;
      put_root_1092 <= 0;
      put_isFree_1093 <= 0;
      put_index_1094 <= 0;
      put_size_1095 <= 0;
      put_isLeaf_1096 <= 0;
      put_nextFree_1097 <= 0;
      put_Key_0_1098 <= 0;
      put_KeyCompares_0_1099 <= 0;
      put_KeyCollapse_0_1100 <= 0;
      put_Data_0_1101 <= 0;
      put_Key_1_1102 <= 0;
      put_KeyCompares_1_1103 <= 0;
      put_KeyCollapse_1_1104 <= 0;
      put_Data_1_1105 <= 0;
      put_Key_2_1106 <= 0;
      put_KeyCompares_2_1107 <= 0;
      put_KeyCollapse_2_1108 <= 0;
      put_Data_2_1109 <= 0;
      put_Key_3_1110 <= 0;
      put_KeyCompares_3_1111 <= 0;
      put_KeyCollapse_3_1112 <= 0;
      put_Data_3_1113 <= 0;
      put_Found_1114 <= 0;
      put_Key_1115 <= 0;
      put_FoundKey_1116 <= 0;
      put_Data_1117 <= 0;
      put_BtreeIndex_1118 <= 0;
      put_StuckIndex_1119 <= 0;
      put_MergeSuccess_1120 <= 0;
      put_index_1121 <= 0;
      put_size_1122 <= 0;
      put_isLeaf_1123 <= 0;
      put_nextFree_1124 <= 0;
      put_Key_0_1125 <= 0;
      put_KeyCompares_0_1126 <= 0;
      put_KeyCollapse_0_1127 <= 0;
      put_Data_0_1128 <= 0;
      put_Key_1_1129 <= 0;
      put_KeyCompares_1_1130 <= 0;
      put_KeyCollapse_1_1131 <= 0;
      put_Data_1_1132 <= 0;
      put_Key_2_1133 <= 0;
      put_KeyCompares_2_1134 <= 0;
      put_KeyCollapse_2_1135 <= 0;
      put_Data_2_1136 <= 0;
      put_Key_3_1137 <= 0;
      put_KeyCompares_3_1138 <= 0;
      put_KeyCollapse_3_1139 <= 0;
      put_Data_3_1140 <= 0;
      put_Found_1141 <= 0;
      put_Key_1142 <= 0;
      put_FoundKey_1143 <= 0;
      put_Data_1144 <= 0;
      put_BtreeIndex_1145 <= 0;
      put_StuckIndex_1146 <= 0;
      put_MergeSuccess_1147 <= 0;
      put_childKey_1148 <= 0;
      put_childData_1149 <= 0;
      put_indexLeft_1150 <= 0;
      put_indexRight_1151 <= 0;
      put_midKey_1152 <= 0;
      put_success_1153 <= 0;
      put_test_1154 <= 0;
      put_next_1155 <= 0;
      put_root_1156 <= 0;
      put_isFree_1157 <= 0;
      put_index_1158 <= 0;
      put_size_1159 <= 0;
      put_isLeaf_1160 <= 0;
      put_nextFree_1161 <= 0;
      put_Key_0_1162 <= 0;
      put_KeyCompares_0_1163 <= 0;
      put_KeyCollapse_0_1164 <= 0;
      put_Data_0_1165 <= 0;
      put_Key_1_1166 <= 0;
      put_KeyCompares_1_1167 <= 0;
      put_KeyCollapse_1_1168 <= 0;
      put_Data_1_1169 <= 0;
      put_Key_2_1170 <= 0;
      put_KeyCompares_2_1171 <= 0;
      put_KeyCollapse_2_1172 <= 0;
      put_Data_2_1173 <= 0;
      put_Key_3_1174 <= 0;
      put_KeyCompares_3_1175 <= 0;
      put_KeyCollapse_3_1176 <= 0;
      put_Data_3_1177 <= 0;
      put_Found_1178 <= 0;
      put_Key_1179 <= 0;
      put_FoundKey_1180 <= 0;
      put_Data_1181 <= 0;
      put_BtreeIndex_1182 <= 0;
      put_StuckIndex_1183 <= 0;
      put_MergeSuccess_1184 <= 0;
      put_index_1185 <= 0;
      put_size_1186 <= 0;
      put_isLeaf_1187 <= 0;
      put_nextFree_1188 <= 0;
      put_Key_0_1189 <= 0;
      put_KeyCompares_0_1190 <= 0;
      put_KeyCollapse_0_1191 <= 0;
      put_Data_0_1192 <= 0;
      put_Key_1_1193 <= 0;
      put_KeyCompares_1_1194 <= 0;
      put_KeyCollapse_1_1195 <= 0;
      put_Data_1_1196 <= 0;
      put_Key_2_1197 <= 0;
      put_KeyCompares_2_1198 <= 0;
      put_KeyCollapse_2_1199 <= 0;
      put_Data_2_1200 <= 0;
      put_Key_3_1201 <= 0;
      put_KeyCompares_3_1202 <= 0;
      put_KeyCollapse_3_1203 <= 0;
      put_Data_3_1204 <= 0;
      put_Found_1205 <= 0;
      put_Key_1206 <= 0;
      put_FoundKey_1207 <= 0;
      put_Data_1208 <= 0;
      put_BtreeIndex_1209 <= 0;
      put_StuckIndex_1210 <= 0;
      put_MergeSuccess_1211 <= 0;
      put_childKey_1212 <= 0;
      put_leftChild_1213 <= 0;
      put_rightChild_1214 <= 0;
      put_childData_1215 <= 0;
      put_indexLeft_1216 <= 0;
      put_indexRight_1217 <= 0;
      put_midKey_1218 <= 0;
      put_success_1219 <= 0;
      put_test_1220 <= 0;
      put_next_1221 <= 0;
      put_root_1222 <= 0;
      put_isFree_1223 <= 0;
      put_index_1224 <= 0;
      put_size_1225 <= 0;
      put_isLeaf_1226 <= 0;
      put_nextFree_1227 <= 0;
      put_Key_0_1228 <= 0;
      put_KeyCompares_0_1229 <= 0;
      put_KeyCollapse_0_1230 <= 0;
      put_Data_0_1231 <= 0;
      put_Key_1_1232 <= 0;
      put_KeyCompares_1_1233 <= 0;
      put_KeyCollapse_1_1234 <= 0;
      put_Data_1_1235 <= 0;
      put_Key_2_1236 <= 0;
      put_KeyCompares_2_1237 <= 0;
      put_KeyCollapse_2_1238 <= 0;
      put_Data_2_1239 <= 0;
      put_Key_3_1240 <= 0;
      put_KeyCompares_3_1241 <= 0;
      put_KeyCollapse_3_1242 <= 0;
      put_Data_3_1243 <= 0;
      put_Found_1244 <= 0;
      put_Key_1245 <= 0;
      put_FoundKey_1246 <= 0;
      put_Data_1247 <= 0;
      put_BtreeIndex_1248 <= 0;
      put_StuckIndex_1249 <= 0;
      put_MergeSuccess_1250 <= 0;
      put_index_1251 <= 0;
      put_size_1252 <= 0;
      put_isLeaf_1253 <= 0;
      put_nextFree_1254 <= 0;
      put_Key_0_1255 <= 0;
      put_KeyCompares_0_1256 <= 0;
      put_KeyCollapse_0_1257 <= 0;
      put_Data_0_1258 <= 0;
      put_Key_1_1259 <= 0;
      put_KeyCompares_1_1260 <= 0;
      put_KeyCollapse_1_1261 <= 0;
      put_Data_1_1262 <= 0;
      put_Key_2_1263 <= 0;
      put_KeyCompares_2_1264 <= 0;
      put_KeyCollapse_2_1265 <= 0;
      put_Data_2_1266 <= 0;
      put_Key_3_1267 <= 0;
      put_KeyCompares_3_1268 <= 0;
      put_KeyCollapse_3_1269 <= 0;
      put_Data_3_1270 <= 0;
      put_Found_1271 <= 0;
      put_Key_1272 <= 0;
      put_FoundKey_1273 <= 0;
      put_Data_1274 <= 0;
      put_BtreeIndex_1275 <= 0;
      put_StuckIndex_1276 <= 0;
      put_MergeSuccess_1277 <= 0;
      put_childKey_1278 <= 0;
      put_childData_1279 <= 0;
      put_indexLeft_1280 <= 0;
      put_indexRight_1281 <= 0;
      put_midKey_1282 <= 0;
      put_success_1283 <= 0;
      put_test_1284 <= 0;
      put_next_1285 <= 0;
      put_root_1286 <= 0;
      put_isFree_1287 <= 0;
      put_index_1288 <= 0;
      put_size_1289 <= 0;
      put_isLeaf_1290 <= 0;
      put_nextFree_1291 <= 0;
      put_Key_0_1292 <= 0;
      put_KeyCompares_0_1293 <= 0;
      put_KeyCollapse_0_1294 <= 0;
      put_Data_0_1295 <= 0;
      put_Key_1_1296 <= 0;
      put_KeyCompares_1_1297 <= 0;
      put_KeyCollapse_1_1298 <= 0;
      put_Data_1_1299 <= 0;
      put_Key_2_1300 <= 0;
      put_KeyCompares_2_1301 <= 0;
      put_KeyCollapse_2_1302 <= 0;
      put_Data_2_1303 <= 0;
      put_Key_3_1304 <= 0;
      put_KeyCompares_3_1305 <= 0;
      put_KeyCollapse_3_1306 <= 0;
      put_Data_3_1307 <= 0;
      put_Found_1308 <= 0;
      put_Key_1309 <= 0;
      put_FoundKey_1310 <= 0;
      put_Data_1311 <= 0;
      put_BtreeIndex_1312 <= 0;
      put_StuckIndex_1313 <= 0;
      put_MergeSuccess_1314 <= 0;
      put_index_1315 <= 0;
      put_size_1316 <= 0;
      put_isLeaf_1317 <= 0;
      put_nextFree_1318 <= 0;
      put_Key_0_1319 <= 0;
      put_KeyCompares_0_1320 <= 0;
      put_KeyCollapse_0_1321 <= 0;
      put_Data_0_1322 <= 0;
      put_Key_1_1323 <= 0;
      put_KeyCompares_1_1324 <= 0;
      put_KeyCollapse_1_1325 <= 0;
      put_Data_1_1326 <= 0;
      put_Key_2_1327 <= 0;
      put_KeyCompares_2_1328 <= 0;
      put_KeyCollapse_2_1329 <= 0;
      put_Data_2_1330 <= 0;
      put_Key_3_1331 <= 0;
      put_KeyCompares_3_1332 <= 0;
      put_KeyCollapse_3_1333 <= 0;
      put_Data_3_1334 <= 0;
      put_Found_1335 <= 0;
      put_Key_1336 <= 0;
      put_FoundKey_1337 <= 0;
      put_Data_1338 <= 0;
      put_BtreeIndex_1339 <= 0;
      put_StuckIndex_1340 <= 0;
      put_MergeSuccess_1341 <= 0;
      put_childKey_1342 <= 0;
      put_leftChild_1343 <= 0;
      put_rightChild_1344 <= 0;
      put_childData_1345 <= 0;
      put_indexLeft_1346 <= 0;
      put_indexRight_1347 <= 0;
      put_midKey_1348 <= 0;
      put_success_1349 <= 0;
      put_test_1350 <= 0;
      put_next_1351 <= 0;
      put_root_1352 <= 0;
      put_isFree_1353 <= 0;
      put_index_1354 <= 0;
      put_size_1355 <= 0;
      put_isLeaf_1356 <= 0;
      put_nextFree_1357 <= 0;
      put_Key_0_1358 <= 0;
      put_KeyCompares_0_1359 <= 0;
      put_KeyCollapse_0_1360 <= 0;
      put_Data_0_1361 <= 0;
      put_Key_1_1362 <= 0;
      put_KeyCompares_1_1363 <= 0;
      put_KeyCollapse_1_1364 <= 0;
      put_Data_1_1365 <= 0;
      put_Key_2_1366 <= 0;
      put_KeyCompares_2_1367 <= 0;
      put_KeyCollapse_2_1368 <= 0;
      put_Data_2_1369 <= 0;
      put_Key_3_1370 <= 0;
      put_KeyCompares_3_1371 <= 0;
      put_KeyCollapse_3_1372 <= 0;
      put_Data_3_1373 <= 0;
      put_Found_1374 <= 0;
      put_Key_1375 <= 0;
      put_FoundKey_1376 <= 0;
      put_Data_1377 <= 0;
      put_BtreeIndex_1378 <= 0;
      put_StuckIndex_1379 <= 0;
      put_MergeSuccess_1380 <= 0;
      put_index_1381 <= 0;
      put_size_1382 <= 0;
      put_isLeaf_1383 <= 0;
      put_nextFree_1384 <= 0;
      put_Key_0_1385 <= 0;
      put_KeyCompares_0_1386 <= 0;
      put_KeyCollapse_0_1387 <= 0;
      put_Data_0_1388 <= 0;
      put_Key_1_1389 <= 0;
      put_KeyCompares_1_1390 <= 0;
      put_KeyCollapse_1_1391 <= 0;
      put_Data_1_1392 <= 0;
      put_Key_2_1393 <= 0;
      put_KeyCompares_2_1394 <= 0;
      put_KeyCollapse_2_1395 <= 0;
      put_Data_2_1396 <= 0;
      put_Key_3_1397 <= 0;
      put_KeyCompares_3_1398 <= 0;
      put_KeyCollapse_3_1399 <= 0;
      put_Data_3_1400 <= 0;
      put_Found_1401 <= 0;
      put_Key_1402 <= 0;
      put_FoundKey_1403 <= 0;
      put_Data_1404 <= 0;
      put_BtreeIndex_1405 <= 0;
      put_StuckIndex_1406 <= 0;
      put_MergeSuccess_1407 <= 0;
      put_childKey_1408 <= 0;
      put_childData_1409 <= 0;
      put_indexLeft_1410 <= 0;
      put_indexRight_1411 <= 0;
      put_midKey_1412 <= 0;
      put_success_1413 <= 0;
      put_test_1414 <= 0;
      put_next_1415 <= 0;
      put_root_1416 <= 0;
      put_isFree_1417 <= 0;
      put_index_1418 <= 0;
      put_size_1419 <= 0;
      put_isLeaf_1420 <= 0;
      put_nextFree_1421 <= 0;
      put_Key_0_1422 <= 0;
      put_KeyCompares_0_1423 <= 0;
      put_KeyCollapse_0_1424 <= 0;
      put_Data_0_1425 <= 0;
      put_Key_1_1426 <= 0;
      put_KeyCompares_1_1427 <= 0;
      put_KeyCollapse_1_1428 <= 0;
      put_Data_1_1429 <= 0;
      put_Key_2_1430 <= 0;
      put_KeyCompares_2_1431 <= 0;
      put_KeyCollapse_2_1432 <= 0;
      put_Data_2_1433 <= 0;
      put_Key_3_1434 <= 0;
      put_KeyCompares_3_1435 <= 0;
      put_KeyCollapse_3_1436 <= 0;
      put_Data_3_1437 <= 0;
      put_Found_1438 <= 0;
      put_Key_1439 <= 0;
      put_FoundKey_1440 <= 0;
      put_Data_1441 <= 0;
      put_BtreeIndex_1442 <= 0;
      put_StuckIndex_1443 <= 0;
      put_MergeSuccess_1444 <= 0;
      put_index_1445 <= 0;
      put_size_1446 <= 0;
      put_isLeaf_1447 <= 0;
      put_nextFree_1448 <= 0;
      put_Key_0_1449 <= 0;
      put_KeyCompares_0_1450 <= 0;
      put_KeyCollapse_0_1451 <= 0;
      put_Data_0_1452 <= 0;
      put_Key_1_1453 <= 0;
      put_KeyCompares_1_1454 <= 0;
      put_KeyCollapse_1_1455 <= 0;
      put_Data_1_1456 <= 0;
      put_Key_2_1457 <= 0;
      put_KeyCompares_2_1458 <= 0;
      put_KeyCollapse_2_1459 <= 0;
      put_Data_2_1460 <= 0;
      put_Key_3_1461 <= 0;
      put_KeyCompares_3_1462 <= 0;
      put_KeyCollapse_3_1463 <= 0;
      put_Data_3_1464 <= 0;
      put_Found_1465 <= 0;
      put_Key_1466 <= 0;
      put_FoundKey_1467 <= 0;
      put_Data_1468 <= 0;
      put_BtreeIndex_1469 <= 0;
      put_StuckIndex_1470 <= 0;
      put_MergeSuccess_1471 <= 0;
      put_childKey_1472 <= 0;
      put_leftChild_1473 <= 0;
      put_rightChild_1474 <= 0;
      put_childData_1475 <= 0;
      put_indexLeft_1476 <= 0;
      put_indexRight_1477 <= 0;
      put_midKey_1478 <= 0;
      put_success_1479 <= 0;
      put_test_1480 <= 0;
      put_next_1481 <= 0;
      put_root_1482 <= 0;
      put_isFree_1483 <= 0;
      stuckIsLeaf_7_requestedAt <= -1;
      stuckIsLeaf_8_requestedAt <= -1;
      stuckIsFree_11_requestedAt <= -1;
      freeNext_9_requestedAt <= -1;
      freeNext_10_requestedAt <= -1;
      stuckSize_5_requestedAt <= -1;
      stuckSize_6_requestedAt <= -1;
      stuckKeys_1_requestedAt <= -1;
      stuckKeys_2_requestedAt <= -1;
      stuckData_3_requestedAt <= -1;
      stuckData_4_requestedAt <= -1;
    end
    else if (processCurrent == 6) begin
      case(put_pc)
        0: begin
          put_k_0 <= put_k_0+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0806:<init>|  Chip.java:0805:Inc|  Btree.java:6068:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        1: begin
          put_d_1 <= put_k_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:6068:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        2: begin
          put_d_1 <= put_d_1+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0806:<init>|  Chip.java:0805:Inc|  Btree.java:6068:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        3: begin
          put_BtreeIndex_100 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2250:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        4: begin
          put_index_76 <= put_BtreeIndex_100;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        5: begin
          put_stuckSize_5_index_36 <= put_index_76;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_76;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_76;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_76;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        6: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        7: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        8: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        9: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        10: begin
          put_size_77 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_78 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_80 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_83 <= stuckData_stuckData_3_result_0;
          put_Key_1_84 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_87 <= stuckData_stuckData_3_result_1;
          put_Key_2_88 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_91 <= stuckData_stuckData_3_result_2;
          put_Key_3_92 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_95 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        11: begin
          if (put_isLeaf_78 == 0) begin
            put_pc <= 18;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        12: begin
          put_KeyCompares_0_81 <= put_k_0 == put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 == put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 == put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 == put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0801:<init>|  Btree.java:0800:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        13: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        14: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        15: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Key_97 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Key_97 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Key_97 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Key_97 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0844:<init>|  Btree.java:0843:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        16: begin
          put_pc <= 24;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2258:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        17: begin
          put_pc <= 24;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        18: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        19: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        20: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        21: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        22: begin
          put_BtreeIndex_100 <= put_Data_99;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2262:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        23: begin
          put_pc <= 4;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2263:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        24: begin
          if (put_Found_96 == 0) begin
            put_pc <= 27;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        25: begin
          if (put_StuckIndex_101 == put_size_77) begin
            put_size_77 <= put_size_77+1;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2293:Then|  Chip.java:0610:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        26: begin
          put_pc <= 38;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        27: begin
          put_notFull_109 <= put_size_77< 4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:2297:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        28: begin
          if (put_notFull_109 == 0) begin
            put_pc <= 37;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        29: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        30: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        31: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        32: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        33: begin
          put_size_77 <= put_size_77+1;
          if (3 > put_StuckIndex_101) begin
            put_Key_3_92 <= put_Key_2_88;
            put_Data_3_95 <= put_Data_2_91;
          end
          if (2 > put_StuckIndex_101) begin
            put_Key_2_88 <= put_Key_1_84;
            put_Data_2_91 <= put_Data_1_87;
          end
          if (1 > put_StuckIndex_101) begin
            put_Key_1_84 <= put_Key_0_80;
            put_Data_1_87 <= put_Data_0_83;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0700:<init>|  Btree.java:0699:InsertElementAt|  Btree.java:2302:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        34: begin
          put_Found_96 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        35: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0592:<init>|  Chip.java:0591:COntinue|  Btree.java:2304:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        36: begin
          put_pc <= 38;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        37: begin
          put_pc <= 42;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2307:Else|  Chip.java:0620:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        38: begin
          put_stuckSize_6_index_37 <= put_index_76;
          put_stuckSize_6_value_38 <= put_size_77;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_76;
          put_stuckKeys_2_value_26 <= put_Key_0_80;
          put_stuckKeys_2_value_27 <= put_Key_1_84;
          put_stuckKeys_2_value_28 <= put_Key_2_88;
          put_stuckKeys_2_value_29 <= put_Key_3_92;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_76;
          put_stuckData_4_value_32 <= put_Data_0_83;
          put_stuckData_4_value_33 <= put_Data_1_87;
          put_stuckData_4_value_34 <= put_Data_2_91;
          put_stuckData_4_value_35 <= put_Data_3_95;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        39: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        40: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        41: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2329:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        42: begin
          if (put_Found_96 >  0) begin
            put_pc <= 450;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0578:<init>|  Chip.java:0577:GONotZero|  Btree.java:2334:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        43: begin
          if (put_BtreeIndex_100 == 0) begin
            put_pc <= 45;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        44: begin
          put_pc <= 138;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        45: begin
          put_index_110 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        46: begin
          put_stuckSize_5_index_36 <= put_index_110;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_110;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_110;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_110;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        47: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        48: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        49: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        50: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        51: begin
          put_size_111 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_112 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_114 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_117 <= stuckData_stuckData_3_result_0;
          put_Key_1_118 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_121 <= stuckData_stuckData_3_result_1;
          put_Key_2_122 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_125 <= stuckData_stuckData_3_result_2;
          put_Key_3_126 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_129 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1525:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        52: begin
          if (put_size_111 < 4) begin
            put_pc <= 98;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1530:<init>|  Btree.java:1529:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        53: begin
          put_Key_0_141 <= put_Key_0_114;
          put_Data_0_144 <= put_Data_0_117;
          put_Key_1_145 <= put_Key_1_118;
          put_Data_1_148 <= put_Data_1_121;
          put_size_138 <= 2;
          put_Key_0_168 <= put_Key_2_122;
          put_Data_0_171 <= put_Data_2_125;
          put_Key_1_172 <= put_Key_3_126;
          put_Data_1_175 <= put_Data_3_129;
          put_size_165 <= 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1041:<init>|  Btree.java:1040:splitIntoTwo|  Btree.java:1547:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        54: begin
          put_root_199 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        55: begin
          put_freeNext_9_index_194 <= put_root_199;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        56: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        57: begin
          put_indexLeft_191 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        58: begin
          if (put_indexLeft_191 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_201 <= 1;
          put_isFree_202 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        59: begin
          put_freeNext_9_index_194 <= put_indexLeft_191;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_191;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_201;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_191;
          put_stuckIsFree_11_value_198 <= put_isFree_202;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        60: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        61: begin
          put_next_200 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        62: begin
          put_freeNext_10_index_195 <= put_root_199;
          put_freeNext_10_value_196 <= put_next_200;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        63: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        64: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        65: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        66: begin
          put_stuckSize_6_index_37 <= put_indexLeft_191;
          put_stuckSize_6_value_38 <= put_size_138;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_191;
          put_stuckKeys_2_value_26 <= put_Key_0_141;
          put_stuckKeys_2_value_27 <= put_Key_1_145;
          put_stuckKeys_2_value_28 <= put_Key_2_149;
          put_stuckKeys_2_value_29 <= put_Key_3_153;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_191;
          put_stuckData_4_value_32 <= put_Data_0_144;
          put_stuckData_4_value_33 <= put_Data_1_148;
          put_stuckData_4_value_34 <= put_Data_2_152;
          put_stuckData_4_value_35 <= put_Data_3_156;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        67: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        68: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        69: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        70: begin
          put_root_203 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        71: begin
          put_freeNext_9_index_194 <= put_root_203;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        72: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        73: begin
          put_indexRight_192 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        74: begin
          if (put_indexRight_192 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_205 <= 1;
          put_isFree_206 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        75: begin
          put_freeNext_9_index_194 <= put_indexRight_192;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexRight_192;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_205;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexRight_192;
          put_stuckIsFree_11_value_198 <= put_isFree_206;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        76: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        77: begin
          put_next_204 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        78: begin
          put_freeNext_10_index_195 <= put_root_203;
          put_freeNext_10_value_196 <= put_next_204;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        79: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        80: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        81: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        82: begin
          put_stuckSize_6_index_37 <= put_indexRight_192;
          put_stuckSize_6_value_38 <= put_size_165;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexRight_192;
          put_stuckKeys_2_value_26 <= put_Key_0_168;
          put_stuckKeys_2_value_27 <= put_Key_1_172;
          put_stuckKeys_2_value_28 <= put_Key_2_176;
          put_stuckKeys_2_value_29 <= put_Key_3_180;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexRight_192;
          put_stuckData_4_value_32 <= put_Data_0_171;
          put_stuckData_4_value_33 <= put_Data_1_175;
          put_stuckData_4_value_34 <= put_Data_2_179;
          put_stuckData_4_value_35 <= put_Data_3_183;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        83: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        84: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        85: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1550:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        86: begin
          case (put_size_138)
            1: begin
              put_Key_158 <= put_Key_0_141;
              put_Data_160 <= put_Data_0_144;
            end
            2: begin
              put_Key_158 <= put_Key_1_145;
              put_Data_160 <= put_Data_1_148;
            end
            3: begin
              put_Key_158 <= put_Key_2_149;
              put_Data_160 <= put_Data_2_152;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0530:<init>|  Btree.java:0529:LastElement|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        87: begin
          put_Key_185 <= put_Key_0_168;
          put_Data_187 <= put_Data_0_171;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0503:<init>|  Btree.java:0502:FirstElement|  Btree.java:1553:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        88: begin
          put_midKey_193 <= (put_Key_158 + put_Key_185) / 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0833:<init>|  Chip.java:0832:Average|  Btree.java:1554:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        89: begin
          put_size_111 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0394:<init>|  Btree.java:0393:Clear|  Btree.java:1555:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        90: begin
          case (put_size_111)
            0: begin
              put_Key_0_114 <= put_midKey_193;
              put_Data_0_117 <= put_indexLeft_191;
            end
            1: begin
              put_Key_1_118 <= put_midKey_193;
              put_Data_1_121 <= put_indexLeft_191;
            end
            2: begin
              put_Key_2_122 <= put_midKey_193;
              put_Data_2_125 <= put_indexLeft_191;
            end
            3: begin
              put_Key_3_126 <= put_midKey_193;
              put_Data_3_129 <= put_indexLeft_191;
            end
          endcase
          put_size_111 <= put_size_111+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0423:<init>|  Btree.java:0422:Push|  Btree.java:1556:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        91: begin
          case (put_size_111)
            0: begin
              put_Key_0_114 <= put_midKey_193;
              put_Data_0_117 <= put_indexRight_192;
            end
            1: begin
              put_Key_1_118 <= put_midKey_193;
              put_Data_1_121 <= put_indexRight_192;
            end
            2: begin
              put_Key_2_122 <= put_midKey_193;
              put_Data_2_125 <= put_indexRight_192;
            end
            3: begin
              put_Key_3_126 <= put_midKey_193;
              put_Data_3_129 <= put_indexRight_192;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0480:<init>|  Btree.java:0479:SetPastLastElement|  Btree.java:1557:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        92: begin
          put_isLeaf_112 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1558:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        93: begin
          put_stuckSize_6_index_37 <= put_index_110;
          put_stuckSize_6_value_38 <= put_size_111;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_index_110;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_112;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_110;
          put_stuckKeys_2_value_26 <= put_Key_0_114;
          put_stuckKeys_2_value_27 <= put_Key_1_118;
          put_stuckKeys_2_value_28 <= put_Key_2_122;
          put_stuckKeys_2_value_29 <= put_Key_3_126;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_110;
          put_stuckData_4_value_32 <= put_Data_0_117;
          put_stuckData_4_value_33 <= put_Data_1_121;
          put_stuckData_4_value_34 <= put_Data_2_125;
          put_stuckData_4_value_35 <= put_Data_3_129;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1559:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        94: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1559:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        95: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1559:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        96: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1559:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        97: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1559:code|  Chip.java:0530:<init>|  Btree.java:1528:<init>|  Btree.java:1527:splitRootLeaf|  Btree.java:2338:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        98: begin
          put_BtreeIndex_100 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2250:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        99: begin
          put_index_76 <= put_BtreeIndex_100;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        100: begin
          put_stuckSize_5_index_36 <= put_index_76;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_76;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_76;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_76;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        101: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        102: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        103: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        104: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        105: begin
          put_size_77 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_78 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_80 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_83 <= stuckData_stuckData_3_result_0;
          put_Key_1_84 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_87 <= stuckData_stuckData_3_result_1;
          put_Key_2_88 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_91 <= stuckData_stuckData_3_result_2;
          put_Key_3_92 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_95 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        106: begin
          if (put_isLeaf_78 == 0) begin
            put_pc <= 113;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        107: begin
          put_KeyCompares_0_81 <= put_k_0 == put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 == put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 == put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 == put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0801:<init>|  Btree.java:0800:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        108: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        109: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        110: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Key_97 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Key_97 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Key_97 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Key_97 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0844:<init>|  Btree.java:0843:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        111: begin
          put_pc <= 119;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2258:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        112: begin
          put_pc <= 119;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        113: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        114: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        115: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        116: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        117: begin
          put_BtreeIndex_100 <= put_Data_99;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2262:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        118: begin
          put_pc <= 99;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2263:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        119: begin
          if (put_Found_96 == 0) begin
            put_pc <= 122;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        120: begin
          if (put_StuckIndex_101 == put_size_77) begin
            put_size_77 <= put_size_77+1;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2293:Then|  Chip.java:0610:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        121: begin
          put_pc <= 133;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        122: begin
          put_notFull_208 <= put_size_77< 4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:2297:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        123: begin
          if (put_notFull_208 == 0) begin
            put_pc <= 132;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        124: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        125: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        126: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        127: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        128: begin
          put_size_77 <= put_size_77+1;
          if (3 > put_StuckIndex_101) begin
            put_Key_3_92 <= put_Key_2_88;
            put_Data_3_95 <= put_Data_2_91;
          end
          if (2 > put_StuckIndex_101) begin
            put_Key_2_88 <= put_Key_1_84;
            put_Data_2_91 <= put_Data_1_87;
          end
          if (1 > put_StuckIndex_101) begin
            put_Key_1_84 <= put_Key_0_80;
            put_Data_1_87 <= put_Data_0_83;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0700:<init>|  Btree.java:0699:InsertElementAt|  Btree.java:2302:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        129: begin
          put_Found_96 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        130: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0592:<init>|  Chip.java:0591:COntinue|  Btree.java:2304:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        131: begin
          put_pc <= 133;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        132: begin
          put_pc <= 137;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2307:Else|  Chip.java:0620:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        133: begin
          put_stuckSize_6_index_37 <= put_index_76;
          put_stuckSize_6_value_38 <= put_size_77;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_76;
          put_stuckKeys_2_value_26 <= put_Key_0_80;
          put_stuckKeys_2_value_27 <= put_Key_1_84;
          put_stuckKeys_2_value_28 <= put_Key_2_88;
          put_stuckKeys_2_value_29 <= put_Key_3_92;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_76;
          put_stuckData_4_value_32 <= put_Data_0_83;
          put_stuckData_4_value_33 <= put_Data_1_87;
          put_stuckData_4_value_34 <= put_Data_2_91;
          put_stuckData_4_value_35 <= put_Data_3_95;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        134: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        135: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        136: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2339:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        137: begin
          put_pc <= 450;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2337:<init>|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        138: begin
          put_index_4 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        139: begin
          put_stuckSize_5_index_36 <= put_index_4;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_4;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_4;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_4;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        140: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        141: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        142: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        143: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        144: begin
          put_size_5 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_6 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_8 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_11 <= stuckData_stuckData_3_result_0;
          put_Key_1_12 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_15 <= stuckData_stuckData_3_result_1;
          put_Key_2_16 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_19 <= stuckData_stuckData_3_result_2;
          put_Key_3_20 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_23 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2344:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        145: begin
          put_full_107 <= put_size_5>=3 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Ge|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        146: begin
          if (put_full_107 == 0) begin
            put_pc <= 198;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        147: begin
          put_index_209 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        148: begin
          put_stuckSize_5_index_36 <= put_index_209;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_209;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_209;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_209;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        149: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        150: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        151: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        152: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        153: begin
          put_size_210 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_211 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_213 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_216 <= stuckData_stuckData_3_result_0;
          put_Key_1_217 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_220 <= stuckData_stuckData_3_result_1;
          put_Key_2_221 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_224 <= stuckData_stuckData_3_result_2;
          put_Key_3_225 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_228 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1573:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        154: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1576:<init>|  Btree.java:1575:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        155: begin
          put_Key_0_240 <= put_Key_0_213;
          put_Data_0_243 <= put_Data_0_216;
          put_size_237 <= 1;
          put_Data_1_247 <= put_Data_1_220;
          put_Key_0_267 <= put_Key_2_221;
          put_Data_0_270 <= put_Data_2_224;
          case (put_size_210)
            0: begin
              put_size_264 <= -2;
              put_Data_1_274 <= put_Data_3_228;
            end
            1: begin
              put_size_264 <= -1;
              put_Data_1_274 <= put_Data_3_228;
            end
            2: begin
              put_size_264 <= 0;
              put_Data_1_274 <= put_Data_3_228;
            end
            3: begin
              put_size_264 <= 1;
              put_Data_1_274 <= put_Data_3_228;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1078:<init>|  Btree.java:1077:splitIntoThree|  Btree.java:1581:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        156: begin
          put_root_293 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        157: begin
          put_freeNext_9_index_194 <= put_root_293;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        158: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        159: begin
          put_indexLeft_290 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        160: begin
          if (put_indexLeft_290 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_295 <= 0;
          put_isFree_296 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        161: begin
          put_freeNext_9_index_194 <= put_indexLeft_290;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_290;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_295;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_290;
          put_stuckIsFree_11_value_198 <= put_isFree_296;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        162: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        163: begin
          put_next_294 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        164: begin
          put_freeNext_10_index_195 <= put_root_293;
          put_freeNext_10_value_196 <= put_next_294;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        165: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        166: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        167: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        168: begin
          put_stuckSize_6_index_37 <= put_indexLeft_290;
          put_stuckSize_6_value_38 <= put_size_237;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_290;
          put_stuckKeys_2_value_26 <= put_Key_0_240;
          put_stuckKeys_2_value_27 <= put_Key_1_244;
          put_stuckKeys_2_value_28 <= put_Key_2_248;
          put_stuckKeys_2_value_29 <= put_Key_3_252;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_290;
          put_stuckData_4_value_32 <= put_Data_0_243;
          put_stuckData_4_value_33 <= put_Data_1_247;
          put_stuckData_4_value_34 <= put_Data_2_251;
          put_stuckData_4_value_35 <= put_Data_3_255;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        169: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        170: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        171: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1582:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        172: begin
          put_root_297 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        173: begin
          put_freeNext_9_index_194 <= put_root_297;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        174: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        175: begin
          put_indexRight_291 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        176: begin
          if (put_indexRight_291 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_299 <= 0;
          put_isFree_300 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        177: begin
          put_freeNext_9_index_194 <= put_indexRight_291;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexRight_291;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_299;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexRight_291;
          put_stuckIsFree_11_value_198 <= put_isFree_300;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        178: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        179: begin
          put_next_298 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        180: begin
          put_freeNext_10_index_195 <= put_root_297;
          put_freeNext_10_value_196 <= put_next_298;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        181: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        182: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        183: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        184: begin
          put_stuckSize_6_index_37 <= put_indexRight_291;
          put_stuckSize_6_value_38 <= put_size_264;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexRight_291;
          put_stuckKeys_2_value_26 <= put_Key_0_267;
          put_stuckKeys_2_value_27 <= put_Key_1_271;
          put_stuckKeys_2_value_28 <= put_Key_2_275;
          put_stuckKeys_2_value_29 <= put_Key_3_279;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexRight_291;
          put_stuckData_4_value_32 <= put_Data_0_270;
          put_stuckData_4_value_33 <= put_Data_1_274;
          put_stuckData_4_value_34 <= put_Data_2_278;
          put_stuckData_4_value_35 <= put_Data_3_282;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        185: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        186: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        187: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1583:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        188: begin
          put_midKey_292 <= put_Key_1_217;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1585:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        189: begin
          put_size_210 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0394:<init>|  Btree.java:0393:Clear|  Btree.java:1586:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        190: begin
          case (put_size_210)
            0: begin
              put_Key_0_213 <= put_midKey_292;
              put_Data_0_216 <= put_indexLeft_290;
            end
            1: begin
              put_Key_1_217 <= put_midKey_292;
              put_Data_1_220 <= put_indexLeft_290;
            end
            2: begin
              put_Key_2_221 <= put_midKey_292;
              put_Data_2_224 <= put_indexLeft_290;
            end
            3: begin
              put_Key_3_225 <= put_midKey_292;
              put_Data_3_228 <= put_indexLeft_290;
            end
          endcase
          put_size_210 <= put_size_210+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0423:<init>|  Btree.java:0422:Push|  Btree.java:1587:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        191: begin
          case (put_size_210)
            0: begin
              put_Key_0_213 <= put_midKey_292;
              put_Data_0_216 <= put_indexRight_291;
            end
            1: begin
              put_Key_1_217 <= put_midKey_292;
              put_Data_1_220 <= put_indexRight_291;
            end
            2: begin
              put_Key_2_221 <= put_midKey_292;
              put_Data_2_224 <= put_indexRight_291;
            end
            3: begin
              put_Key_3_225 <= put_midKey_292;
              put_Data_3_228 <= put_indexRight_291;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0480:<init>|  Btree.java:0479:SetPastLastElement|  Btree.java:1588:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        192: begin
          put_stuckSize_6_index_37 <= put_index_209;
          put_stuckSize_6_value_38 <= put_size_210;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_209;
          put_stuckKeys_2_value_26 <= put_Key_0_213;
          put_stuckKeys_2_value_27 <= put_Key_1_217;
          put_stuckKeys_2_value_28 <= put_Key_2_221;
          put_stuckKeys_2_value_29 <= put_Key_3_225;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_209;
          put_stuckData_4_value_32 <= put_Data_0_216;
          put_stuckData_4_value_33 <= put_Data_1_220;
          put_stuckData_4_value_34 <= put_Data_2_224;
          put_stuckData_4_value_35 <= put_Data_3_228;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1589:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        193: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1589:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        194: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1589:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        195: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1589:splitRootBranch|  Btree.java:2350:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        196: begin
          put_pc <= 42;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2351:Then|  Chip.java:0610:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        197: begin
          put_pc <= 198;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2349:<init>|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        198: begin
          put_parent_104 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2355:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        199: begin
          put_index_4 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        200: begin
          put_stuckSize_5_index_36 <= put_index_4;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_4;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_4;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_4;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        201: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        202: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        203: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        204: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        205: begin
          put_size_5 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_6 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_8 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_11 <= stuckData_stuckData_3_result_0;
          put_Key_1_12 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_15 <= stuckData_stuckData_3_result_1;
          put_Key_2_16 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_19 <= stuckData_stuckData_3_result_2;
          put_Key_3_20 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_23 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2360:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        206: begin
          put_KeyCompares_0_9 <= put_k_0 <= put_Key_0_8 && 0 < put_size_5;
          put_KeyCollapse_0_10 <= 0;
          put_KeyCompares_1_13 <= put_k_0 >  put_Key_0_8 && put_k_0 <= put_Key_1_12 && 1 < put_size_5;
          put_KeyCollapse_1_14 <= 1;
          put_KeyCompares_2_17 <= put_k_0 >  put_Key_1_12 && put_k_0 <= put_Key_2_16 && 2 < put_size_5;
          put_KeyCollapse_2_18 <= 2;
          put_KeyCompares_3_21 <= put_k_0 >  put_Key_2_16 && put_k_0 <= put_Key_3_20 && 3 < put_size_5;
          put_KeyCollapse_3_22 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2361:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        207: begin
          if (put_KeyCompares_1_13) begin
            put_KeyCompares_0_9 <= 1;
            put_KeyCollapse_0_10 <= put_KeyCollapse_1_14;
          end
          if (put_KeyCompares_3_21) begin
            put_KeyCompares_2_17 <= 1;
            put_KeyCollapse_2_18 <= put_KeyCollapse_3_22;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2361:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        208: begin
          if (put_KeyCompares_2_17) begin
            put_KeyCompares_0_9 <= 1;
            put_KeyCollapse_0_10 <= put_KeyCollapse_2_18;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2361:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        209: begin
          if (put_KeyCompares_0_9) begin
            put_Found_42 <= 1;
            case (put_KeyCollapse_0_10)
              0: begin
                put_StuckIndex_47 <= 0;
                put_FoundKey_44 <= put_Key_0_8;
                put_Data_45 <= put_Data_0_11;
              end
              1: begin
                put_StuckIndex_47 <= 1;
                put_FoundKey_44 <= put_Key_1_12;
                put_Data_45 <= put_Data_1_15;
              end
              2: begin
                put_StuckIndex_47 <= 2;
                put_FoundKey_44 <= put_Key_2_16;
                put_Data_45 <= put_Data_2_19;
              end
              3: begin
                put_StuckIndex_47 <= 3;
                put_FoundKey_44 <= put_Key_3_20;
                put_Data_45 <= put_Data_3_23;
              end
            endcase
          end
          else begin
            put_Found_42 <= 0;
            case (put_size_5)
              0: begin
                put_StuckIndex_47 <= 0;
                put_Data_45 <= put_Data_0_11;
              end
              1: begin
                put_StuckIndex_47 <= 1;
                put_Data_45 <= put_Data_1_15;
              end
              2: begin
                put_StuckIndex_47 <= 2;
                put_Data_45 <= put_Data_2_19;
              end
              3: begin
                put_StuckIndex_47 <= 3;
                put_Data_45 <= put_Data_3_23;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2361:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        210: begin
          put_child_103 <= put_Data_45;
          put_childInparent_105 <= put_StuckIndex_47;
          put_found_106 <= put_Found_42;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2363:<init>|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        211: begin
          put_index_49 <= put_child_103;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        212: begin
          put_stuckSize_5_index_36 <= put_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        213: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        214: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        215: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        216: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        217: begin
          put_size_50 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_56 <= stuckData_stuckData_3_result_0;
          put_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_60 <= stuckData_stuckData_3_result_1;
          put_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_64 <= stuckData_stuckData_3_result_2;
          put_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_68 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2371:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        218: begin
          if (put_isLeaf_51 == 0) begin
            put_pc <= 357;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        219: begin
          put_full_107 <= put_size_50>=4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Ge|  Btree.java:2375:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        220: begin
          if (put_full_107 == 0) begin
            put_pc <= 316;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        221: begin
          if (put_found_106 == 0) begin
            put_pc <= 268;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        222: begin
          put_index_301 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        223: begin
          put_stuckSize_5_index_36 <= put_index_301;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_301;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_301;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_301;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        224: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        225: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        226: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        227: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        228: begin
          put_size_302 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_303 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_305 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_308 <= stuckData_stuckData_3_result_0;
          put_Key_1_309 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_312 <= stuckData_stuckData_3_result_1;
          put_Key_2_313 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_316 <= stuckData_stuckData_3_result_2;
          put_Key_3_317 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_320 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1605:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        229: begin
          case (put_childInparent_105)
            0: begin
              put_childKey_409 <= put_Key_0_305;
              put_childData_410 <= put_Data_0_308;
            end
            1: begin
              put_childKey_409 <= put_Key_1_309;
              put_childData_410 <= put_Data_1_312;
            end
            2: begin
              put_childKey_409 <= put_Key_2_313;
              put_childData_410 <= put_Data_2_316;
            end
            3: begin
              put_childKey_409 <= put_Key_3_317;
              put_childData_410 <= put_Data_3_320;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1608:<init>|  Btree.java:1607:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        230: begin
          put_index_328 <= put_childData_410;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        231: begin
          put_stuckSize_5_index_36 <= put_index_328;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_328;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_328;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_328;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        232: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        233: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        234: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        235: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        236: begin
          put_size_329 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_330 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_332 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_335 <= stuckData_stuckData_3_result_0;
          put_Key_1_336 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_339 <= stuckData_stuckData_3_result_1;
          put_Key_2_340 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_343 <= stuckData_stuckData_3_result_2;
          put_Key_3_344 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_347 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1621:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        237: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1624:<init>|  Btree.java:1623:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        238: begin
          put_Key_0_359 <= put_Key_0_332;
          put_Data_0_362 <= put_Data_0_335;
          put_Key_1_363 <= put_Key_1_336;
          put_Data_1_366 <= put_Data_1_339;
          put_size_356 <= 2;
          put_Key_0_332 <= put_Key_2_340;
          put_Data_0_335 <= put_Data_2_343;
          put_Key_1_336 <= put_Key_3_344;
          put_Data_1_339 <= put_Data_3_347;
          put_size_329 <= 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1124:<init>|  Btree.java:1123:splitLow|  Btree.java:1632:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        239: begin
          put_root_414 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        240: begin
          put_freeNext_9_index_194 <= put_root_414;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        241: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        242: begin
          put_indexLeft_411 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        243: begin
          if (put_indexLeft_411 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_416 <= 1;
          put_isFree_417 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        244: begin
          put_freeNext_9_index_194 <= put_indexLeft_411;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_411;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_416;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_411;
          put_stuckIsFree_11_value_198 <= put_isFree_417;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        245: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        246: begin
          put_next_415 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        247: begin
          put_freeNext_10_index_195 <= put_root_414;
          put_freeNext_10_value_196 <= put_next_415;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        248: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        249: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        250: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        251: begin
          put_stuckSize_6_index_37 <= put_childData_410;
          put_stuckSize_6_value_38 <= put_size_329;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childData_410;
          put_stuckKeys_2_value_26 <= put_Key_0_332;
          put_stuckKeys_2_value_27 <= put_Key_1_336;
          put_stuckKeys_2_value_28 <= put_Key_2_340;
          put_stuckKeys_2_value_29 <= put_Key_3_344;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childData_410;
          put_stuckData_4_value_32 <= put_Data_0_335;
          put_stuckData_4_value_33 <= put_Data_1_339;
          put_stuckData_4_value_34 <= put_Data_2_343;
          put_stuckData_4_value_35 <= put_Data_3_347;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        252: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        253: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        254: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1633:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        255: begin
          put_stuckSize_6_index_37 <= put_indexLeft_411;
          put_stuckSize_6_value_38 <= put_size_356;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_411;
          put_stuckKeys_2_value_26 <= put_Key_0_359;
          put_stuckKeys_2_value_27 <= put_Key_1_363;
          put_stuckKeys_2_value_28 <= put_Key_2_367;
          put_stuckKeys_2_value_29 <= put_Key_3_371;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_411;
          put_stuckData_4_value_32 <= put_Data_0_362;
          put_stuckData_4_value_33 <= put_Data_1_366;
          put_stuckData_4_value_34 <= put_Data_2_370;
          put_stuckData_4_value_35 <= put_Data_3_374;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1634:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        256: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1634:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        257: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1634:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        258: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1634:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        259: begin
          case (put_size_356)
            1: begin
              put_Key_376 <= put_Key_0_359;
              put_Data_378 <= put_Data_0_362;
            end
            2: begin
              put_Key_376 <= put_Key_1_363;
              put_Data_378 <= put_Data_1_366;
            end
            3: begin
              put_Key_376 <= put_Key_2_367;
              put_Data_378 <= put_Data_2_370;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0530:<init>|  Btree.java:0529:LastElement|  Btree.java:1636:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        260: begin
          put_Key_349 <= put_Key_0_332;
          put_Data_351 <= put_Data_0_335;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0503:<init>|  Btree.java:0502:FirstElement|  Btree.java:1637:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        261: begin
          put_midKey_413 <= (put_Key_376 + put_Key_349) / 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0833:<init>|  Chip.java:0832:Average|  Btree.java:1638:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        262: begin
          put_size_302 <= put_size_302+1;
          if (3 > put_childInparent_105) begin
            put_Key_3_317 <= put_Key_2_313;
            put_Data_3_320 <= put_Data_2_316;
          end
          if (2 > put_childInparent_105) begin
            put_Key_2_313 <= put_Key_1_309;
            put_Data_2_316 <= put_Data_1_312;
          end
          if (1 > put_childInparent_105) begin
            put_Key_1_309 <= put_Key_0_305;
            put_Data_1_312 <= put_Data_0_308;
          end
          case (put_childInparent_105)
            0: begin
              put_Key_0_305 <= put_midKey_413;
              put_Data_0_308 <= put_indexLeft_411;
            end
            1: begin
              put_Key_1_309 <= put_midKey_413;
              put_Data_1_312 <= put_indexLeft_411;
            end
            2: begin
              put_Key_2_313 <= put_midKey_413;
              put_Data_2_316 <= put_indexLeft_411;
            end
            3: begin
              put_Key_3_317 <= put_midKey_413;
              put_Data_3_320 <= put_indexLeft_411;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0700:<init>|  Btree.java:0699:InsertElementAt|  Btree.java:1639:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        263: begin
          put_stuckSize_6_index_37 <= put_index_301;
          put_stuckSize_6_value_38 <= put_size_302;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_301;
          put_stuckKeys_2_value_26 <= put_Key_0_305;
          put_stuckKeys_2_value_27 <= put_Key_1_309;
          put_stuckKeys_2_value_28 <= put_Key_2_313;
          put_stuckKeys_2_value_29 <= put_Key_3_317;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_301;
          put_stuckData_4_value_32 <= put_Data_0_308;
          put_stuckData_4_value_33 <= put_Data_1_312;
          put_stuckData_4_value_34 <= put_Data_2_316;
          put_stuckData_4_value_35 <= put_Data_3_320;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1640:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        264: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1640:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        265: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1640:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        266: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1640:splitLeafNotTop|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        267: begin
          put_pc <= 315;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        268: begin
          put_index_418 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        269: begin
          put_stuckSize_5_index_36 <= put_index_418;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_418;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_418;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_418;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        270: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        271: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        272: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        273: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        274: begin
          put_size_419 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_420 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_422 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_425 <= stuckData_stuckData_3_result_0;
          put_Key_1_426 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_429 <= stuckData_stuckData_3_result_1;
          put_Key_2_430 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_433 <= stuckData_stuckData_3_result_2;
          put_Key_3_434 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_437 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1652:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        275: begin
          case (put_size_419)
            0: begin
              put_Key_439 <= put_Key_0_422;
              put_Data_441 <= put_Data_0_425;
            end
            1: begin
              put_Key_439 <= put_Key_1_426;
              put_Data_441 <= put_Data_1_429;
            end
            2: begin
              put_Key_439 <= put_Key_2_430;
              put_Data_441 <= put_Data_2_433;
            end
            3: begin
              put_Key_439 <= put_Key_3_434;
              put_Data_441 <= put_Data_3_437;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0557:<init>|  Btree.java:0556:PastLastElement|  Btree.java:1653:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        276: begin
          put_childIndex_499 <= put_Data_441;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1654:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        277: begin
          put_index_445 <= put_childIndex_499;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        278: begin
          put_stuckSize_5_index_36 <= put_index_445;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_445;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_445;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_445;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        279: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        280: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        281: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        282: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        283: begin
          put_size_446 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_447 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_449 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_452 <= stuckData_stuckData_3_result_0;
          put_Key_1_453 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_456 <= stuckData_stuckData_3_result_1;
          put_Key_2_457 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_460 <= stuckData_stuckData_3_result_2;
          put_Key_3_461 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_464 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1655:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        284: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1658:<init>|  Btree.java:1657:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        285: begin
          put_Key_0_476 <= put_Key_0_449;
          put_Data_0_479 <= put_Data_0_452;
          put_Key_1_480 <= put_Key_1_453;
          put_Data_1_483 <= put_Data_1_456;
          put_size_473 <= 2;
          put_Key_0_449 <= put_Key_2_457;
          put_Data_0_452 <= put_Data_2_460;
          put_Key_1_453 <= put_Key_3_461;
          put_Data_1_456 <= put_Data_3_464;
          put_size_446 <= 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1124:<init>|  Btree.java:1123:splitLow|  Btree.java:1667:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        286: begin
          put_root_502 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        287: begin
          put_freeNext_9_index_194 <= put_root_502;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        288: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        289: begin
          put_leftIndex_500 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        290: begin
          if (put_leftIndex_500 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_504 <= 1;
          put_isFree_505 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        291: begin
          put_freeNext_9_index_194 <= put_leftIndex_500;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_leftIndex_500;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_504;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_leftIndex_500;
          put_stuckIsFree_11_value_198 <= put_isFree_505;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        292: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        293: begin
          put_next_503 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        294: begin
          put_freeNext_10_index_195 <= put_root_502;
          put_freeNext_10_value_196 <= put_next_503;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        295: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        296: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        297: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        298: begin
          put_stuckSize_6_index_37 <= put_leftIndex_500;
          put_stuckSize_6_value_38 <= put_size_473;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_leftIndex_500;
          put_stuckKeys_2_value_26 <= put_Key_0_476;
          put_stuckKeys_2_value_27 <= put_Key_1_480;
          put_stuckKeys_2_value_28 <= put_Key_2_484;
          put_stuckKeys_2_value_29 <= put_Key_3_488;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_leftIndex_500;
          put_stuckData_4_value_32 <= put_Data_0_479;
          put_stuckData_4_value_33 <= put_Data_1_483;
          put_stuckData_4_value_34 <= put_Data_2_487;
          put_stuckData_4_value_35 <= put_Data_3_491;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        299: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        300: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        301: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        302: begin
          put_stuckSize_6_index_37 <= put_childIndex_499;
          put_stuckSize_6_value_38 <= put_size_446;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childIndex_499;
          put_stuckKeys_2_value_26 <= put_Key_0_449;
          put_stuckKeys_2_value_27 <= put_Key_1_453;
          put_stuckKeys_2_value_28 <= put_Key_2_457;
          put_stuckKeys_2_value_29 <= put_Key_3_461;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childIndex_499;
          put_stuckData_4_value_32 <= put_Data_0_452;
          put_stuckData_4_value_33 <= put_Data_1_456;
          put_stuckData_4_value_34 <= put_Data_2_460;
          put_stuckData_4_value_35 <= put_Data_3_464;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        303: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        304: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        305: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1668:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        306: begin
          case (put_size_473)
            1: begin
              put_Key_493 <= put_Key_0_476;
              put_Data_495 <= put_Data_0_479;
            end
            2: begin
              put_Key_493 <= put_Key_1_480;
              put_Data_495 <= put_Data_1_483;
            end
            3: begin
              put_Key_493 <= put_Key_2_484;
              put_Data_495 <= put_Data_2_487;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0530:<init>|  Btree.java:0529:LastElement|  Btree.java:1670:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        307: begin
          put_Key_466 <= put_Key_0_449;
          put_Data_468 <= put_Data_0_452;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0503:<init>|  Btree.java:0502:FirstElement|  Btree.java:1671:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        308: begin
          put_midKey_501 <= (put_Key_493 + put_Key_466) / 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0833:<init>|  Chip.java:0832:Average|  Btree.java:1672:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        309: begin
          case (put_size_419)
            0: begin
              put_Key_0_422 <= put_midKey_501;
              put_Data_0_425 <= put_leftIndex_500;
            end
            1: begin
              put_Key_1_426 <= put_midKey_501;
              put_Data_1_429 <= put_leftIndex_500;
            end
            2: begin
              put_Key_2_430 <= put_midKey_501;
              put_Data_2_433 <= put_leftIndex_500;
            end
            3: begin
              put_Key_3_434 <= put_midKey_501;
              put_Data_3_437 <= put_leftIndex_500;
            end
          endcase
          put_size_419 <= put_size_419+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0423:<init>|  Btree.java:0422:Push|  Btree.java:1673:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        310: begin
          case (put_size_419)
            0: begin
              put_Key_0_422 <= put_midKey_501;
              put_Data_0_425 <= put_childIndex_499;
            end
            1: begin
              put_Key_1_426 <= put_midKey_501;
              put_Data_1_429 <= put_childIndex_499;
            end
            2: begin
              put_Key_2_430 <= put_midKey_501;
              put_Data_2_433 <= put_childIndex_499;
            end
            3: begin
              put_Key_3_434 <= put_midKey_501;
              put_Data_3_437 <= put_childIndex_499;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0480:<init>|  Btree.java:0479:SetPastLastElement|  Btree.java:1674:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        311: begin
          put_stuckSize_6_index_37 <= put_index_418;
          put_stuckSize_6_value_38 <= put_size_419;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_418;
          put_stuckKeys_2_value_26 <= put_Key_0_422;
          put_stuckKeys_2_value_27 <= put_Key_1_426;
          put_stuckKeys_2_value_28 <= put_Key_2_430;
          put_stuckKeys_2_value_29 <= put_Key_3_434;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_418;
          put_stuckData_4_value_32 <= put_Data_0_425;
          put_stuckData_4_value_33 <= put_Data_1_429;
          put_stuckData_4_value_34 <= put_Data_2_433;
          put_stuckData_4_value_35 <= put_Data_3_437;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1675:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        312: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1675:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        313: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1675:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        314: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1675:splitLeafAtTop|  Btree.java:2384:Else|  Chip.java:0620:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Then|  Chip.java:0610:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        315: begin
          put_pc <= 316;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2378:<init>|  Btree.java:2377:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        316: begin
          put_BtreeIndex_100 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2250:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        317: begin
          put_index_76 <= put_BtreeIndex_100;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        318: begin
          put_stuckSize_5_index_36 <= put_index_76;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_76;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_76;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_76;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        319: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        320: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        321: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        322: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        323: begin
          put_size_77 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_78 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_80 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_83 <= stuckData_stuckData_3_result_0;
          put_Key_1_84 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_87 <= stuckData_stuckData_3_result_1;
          put_Key_2_88 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_91 <= stuckData_stuckData_3_result_2;
          put_Key_3_92 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_95 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2254:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        324: begin
          if (put_isLeaf_78 == 0) begin
            put_pc <= 331;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        325: begin
          put_KeyCompares_0_81 <= put_k_0 == put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 == put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 == put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 == put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0801:<init>|  Btree.java:0800:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        326: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        327: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0822:<init>|  Btree.java:0821:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        328: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Key_97 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Key_97 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Key_97 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Key_97 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0844:<init>|  Btree.java:0843:search_eq_parallel|  Btree.java:2257:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        329: begin
          put_pc <= 337;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2258:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        330: begin
          put_pc <= 337;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        331: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        332: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        333: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        334: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2261:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        335: begin
          put_BtreeIndex_100 <= put_Data_99;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2262:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        336: begin
          put_pc <= 317;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2263:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2256:<init>|  Btree.java:2255:code|  Chip.java:0530:<init>|  Btree.java:2253:<init>|  Btree.java:2252:findSearch|  Btree.java:2289:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        337: begin
          if (put_Found_96 == 0) begin
            put_pc <= 340;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        338: begin
          if (put_StuckIndex_101 == put_size_77) begin
            put_size_77 <= put_size_77+1;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2293:Then|  Chip.java:0610:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        339: begin
          put_pc <= 351;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        340: begin
          put_notFull_507 <= put_size_77< 4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:2297:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        341: begin
          if (put_notFull_507 == 0) begin
            put_pc <= 350;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        342: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        343: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        344: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        345: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2301:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        346: begin
          put_size_77 <= put_size_77+1;
          if (3 > put_StuckIndex_101) begin
            put_Key_3_92 <= put_Key_2_88;
            put_Data_3_95 <= put_Data_2_91;
          end
          if (2 > put_StuckIndex_101) begin
            put_Key_2_88 <= put_Key_1_84;
            put_Data_2_91 <= put_Data_1_87;
          end
          if (1 > put_StuckIndex_101) begin
            put_Key_1_84 <= put_Key_0_80;
            put_Data_1_87 <= put_Data_0_83;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0700:<init>|  Btree.java:0699:InsertElementAt|  Btree.java:2302:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        347: begin
          put_Found_96 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        348: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0592:<init>|  Chip.java:0591:COntinue|  Btree.java:2304:Then|  Chip.java:0610:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        349: begin
          put_pc <= 351;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        350: begin
          put_pc <= 355;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2307:Else|  Chip.java:0620:<init>|  Btree.java:2300:<init>|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2292:<init>|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        351: begin
          put_stuckSize_6_index_37 <= put_index_76;
          put_stuckSize_6_value_38 <= put_size_77;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_76;
          put_stuckKeys_2_value_26 <= put_Key_0_80;
          put_stuckKeys_2_value_27 <= put_Key_1_84;
          put_stuckKeys_2_value_28 <= put_Key_2_88;
          put_stuckKeys_2_value_29 <= put_Key_3_92;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_76;
          put_stuckData_4_value_32 <= put_Data_0_83;
          put_stuckData_4_value_33 <= put_Data_1_87;
          put_stuckData_4_value_34 <= put_Data_2_91;
          put_stuckData_4_value_35 <= put_Data_3_95;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        352: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        353: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        354: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:2312:code|  Chip.java:0530:<init>|  Btree.java:2288:<init>|  Btree.java:2287:findAndInsert|  Btree.java:2389:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        355: begin
          put_pc <= 450;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2390:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        356: begin
          put_pc <= 450;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        357: begin
          put_full_107 <= put_size_50>=3 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Ge|  Btree.java:2394:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        358: begin
          if (put_full_107 == 0) begin
            put_pc <= 448;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        359: begin
          if (put_found_106 == 0) begin
            put_pc <= 403;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        360: begin
          put_index_508 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        361: begin
          put_stuckSize_5_index_36 <= put_index_508;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_508;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_508;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_508;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        362: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        363: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        364: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        365: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        366: begin
          put_size_509 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_510 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_512 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_515 <= stuckData_stuckData_3_result_0;
          put_Key_1_516 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_519 <= stuckData_stuckData_3_result_1;
          put_Key_2_520 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_523 <= stuckData_stuckData_3_result_2;
          put_Key_3_524 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_527 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1691:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        367: begin
          case (put_childInparent_105)
            0: begin
              put_childKey_616 <= put_Key_0_512;
              put_childData_617 <= put_Data_0_515;
            end
            1: begin
              put_childKey_616 <= put_Key_1_516;
              put_childData_617 <= put_Data_1_519;
            end
            2: begin
              put_childKey_616 <= put_Key_2_520;
              put_childData_617 <= put_Data_2_523;
            end
            3: begin
              put_childKey_616 <= put_Key_3_524;
              put_childData_617 <= put_Data_3_527;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1693:<init>|  Btree.java:1692:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        368: begin
          put_index_535 <= put_childData_617;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        369: begin
          put_stuckSize_5_index_36 <= put_index_535;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_535;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_535;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_535;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        370: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        371: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        372: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        373: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        374: begin
          put_size_536 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_537 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_539 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_542 <= stuckData_stuckData_3_result_0;
          put_Key_1_543 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_546 <= stuckData_stuckData_3_result_1;
          put_Key_2_547 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_550 <= stuckData_stuckData_3_result_2;
          put_Key_3_551 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_554 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1706:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        375: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1709:<init>|  Btree.java:1708:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        376: begin
          put_Key_0_566 <= put_Key_0_539;
          put_Data_0_569 <= put_Data_0_542;
          put_size_563 <= 1;
          put_Data_1_573 <= put_Data_1_546;
          put_childKey_616 <= put_Key_1_543;
          put_Key_0_539 <= put_Key_2_547;
          put_Data_0_542 <= put_Data_2_550;
          put_Key_1_543 <= put_Key_3_551;
          put_Data_1_546 <= put_Data_3_554;
          put_size_536 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1165:<init>|  Btree.java:1164:splitLowButOne|  Btree.java:1718:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        377: begin
          put_root_621 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        378: begin
          put_freeNext_9_index_194 <= put_root_621;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        379: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        380: begin
          put_indexLeft_618 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        381: begin
          if (put_indexLeft_618 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_623 <= 0;
          put_isFree_624 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        382: begin
          put_freeNext_9_index_194 <= put_indexLeft_618;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_618;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_623;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_618;
          put_stuckIsFree_11_value_198 <= put_isFree_624;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        383: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        384: begin
          put_next_622 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        385: begin
          put_freeNext_10_index_195 <= put_root_621;
          put_freeNext_10_value_196 <= put_next_622;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        386: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        387: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        388: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        389: begin
          put_stuckSize_6_index_37 <= put_indexLeft_618;
          put_stuckSize_6_value_38 <= put_size_563;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_618;
          put_stuckKeys_2_value_26 <= put_Key_0_566;
          put_stuckKeys_2_value_27 <= put_Key_1_570;
          put_stuckKeys_2_value_28 <= put_Key_2_574;
          put_stuckKeys_2_value_29 <= put_Key_3_578;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_618;
          put_stuckData_4_value_32 <= put_Data_0_569;
          put_stuckData_4_value_33 <= put_Data_1_573;
          put_stuckData_4_value_34 <= put_Data_2_577;
          put_stuckData_4_value_35 <= put_Data_3_581;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        390: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        391: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        392: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1719:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        393: begin
          put_stuckSize_6_index_37 <= put_childData_617;
          put_stuckSize_6_value_38 <= put_size_536;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childData_617;
          put_stuckKeys_2_value_26 <= put_Key_0_539;
          put_stuckKeys_2_value_27 <= put_Key_1_543;
          put_stuckKeys_2_value_28 <= put_Key_2_547;
          put_stuckKeys_2_value_29 <= put_Key_3_551;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childData_617;
          put_stuckData_4_value_32 <= put_Data_0_542;
          put_stuckData_4_value_33 <= put_Data_1_546;
          put_stuckData_4_value_34 <= put_Data_2_550;
          put_stuckData_4_value_35 <= put_Data_3_554;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1720:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        394: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1720:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        395: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1720:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        396: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1720:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        397: begin
          put_size_509 <= put_size_509+1;
          if (3 > put_childInparent_105) begin
            put_Key_3_524 <= put_Key_2_520;
            put_Data_3_527 <= put_Data_2_523;
          end
          if (2 > put_childInparent_105) begin
            put_Key_2_520 <= put_Key_1_516;
            put_Data_2_523 <= put_Data_1_519;
          end
          if (1 > put_childInparent_105) begin
            put_Key_1_516 <= put_Key_0_512;
            put_Data_1_519 <= put_Data_0_515;
          end
          case (put_childInparent_105)
            0: begin
              put_Key_0_512 <= put_childKey_616;
              put_Data_0_515 <= put_indexLeft_618;
            end
            1: begin
              put_Key_1_516 <= put_childKey_616;
              put_Data_1_519 <= put_indexLeft_618;
            end
            2: begin
              put_Key_2_520 <= put_childKey_616;
              put_Data_2_523 <= put_indexLeft_618;
            end
            3: begin
              put_Key_3_524 <= put_childKey_616;
              put_Data_3_527 <= put_indexLeft_618;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0700:<init>|  Btree.java:0699:InsertElementAt|  Btree.java:1722:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        398: begin
          put_stuckSize_6_index_37 <= put_index_508;
          put_stuckSize_6_value_38 <= put_size_509;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_508;
          put_stuckKeys_2_value_26 <= put_Key_0_512;
          put_stuckKeys_2_value_27 <= put_Key_1_516;
          put_stuckKeys_2_value_28 <= put_Key_2_520;
          put_stuckKeys_2_value_29 <= put_Key_3_524;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_508;
          put_stuckData_4_value_32 <= put_Data_0_515;
          put_stuckData_4_value_33 <= put_Data_1_519;
          put_stuckData_4_value_34 <= put_Data_2_523;
          put_stuckData_4_value_35 <= put_Data_3_527;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1723:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        399: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1723:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        400: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1723:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        401: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1723:splitBranchNotTop|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        402: begin
          put_pc <= 447;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        403: begin
          put_index_625 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        404: begin
          put_stuckSize_5_index_36 <= put_index_625;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_625;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_625;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_625;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        405: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        406: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        407: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        408: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        409: begin
          put_size_626 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_627 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_629 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_632 <= stuckData_stuckData_3_result_0;
          put_Key_1_633 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_636 <= stuckData_stuckData_3_result_1;
          put_Key_2_637 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_640 <= stuckData_stuckData_3_result_2;
          put_Key_3_641 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_644 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1738:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        410: begin
          case (put_size_626)
            0: begin
              put_Key_646 <= put_Key_0_629;
              put_Data_648 <= put_Data_0_632;
            end
            1: begin
              put_Key_646 <= put_Key_1_633;
              put_Data_648 <= put_Data_1_636;
            end
            2: begin
              put_Key_646 <= put_Key_2_637;
              put_Data_648 <= put_Data_2_640;
            end
            3: begin
              put_Key_646 <= put_Key_3_641;
              put_Data_648 <= put_Data_3_644;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0557:<init>|  Btree.java:0556:PastLastElement|  Btree.java:1740:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        411: begin
          put_childData_734 <= put_Data_648;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1741:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        412: begin
          put_index_652 <= put_childData_734;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        413: begin
          put_stuckSize_5_index_36 <= put_index_652;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_652;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_652;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_652;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        414: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        415: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        416: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        417: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        418: begin
          put_size_653 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_654 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_656 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_659 <= stuckData_stuckData_3_result_0;
          put_Key_1_660 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_663 <= stuckData_stuckData_3_result_1;
          put_Key_2_664 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_667 <= stuckData_stuckData_3_result_2;
          put_Key_3_668 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_671 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1742:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        419: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1745:<init>|  Btree.java:1744:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        420: begin
          put_Key_0_683 <= put_Key_0_656;
          put_Data_0_686 <= put_Data_0_659;
          put_size_680 <= 1;
          put_Data_1_690 <= put_Data_1_663;
          put_midKey_737 <= put_Key_1_660;
          put_Key_0_656 <= put_Key_2_664;
          put_Data_0_659 <= put_Data_2_667;
          put_Key_1_660 <= put_Key_3_668;
          put_Data_1_663 <= put_Data_3_671;
          put_size_653 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1165:<init>|  Btree.java:1164:splitLowButOne|  Btree.java:1754:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        421: begin
          put_root_738 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        422: begin
          put_freeNext_9_index_194 <= put_root_738;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        423: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        424: begin
          put_indexLeft_735 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        425: begin
          if (put_indexLeft_735 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_740 <= 0;
          put_isFree_741 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        426: begin
          put_freeNext_9_index_194 <= put_indexLeft_735;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_735;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_740;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_735;
          put_stuckIsFree_11_value_198 <= put_isFree_741;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        427: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        428: begin
          put_next_739 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        429: begin
          put_freeNext_10_index_195 <= put_root_738;
          put_freeNext_10_value_196 <= put_next_739;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        430: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        431: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        432: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        433: begin
          put_stuckSize_6_index_37 <= put_indexLeft_735;
          put_stuckSize_6_value_38 <= put_size_680;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_735;
          put_stuckKeys_2_value_26 <= put_Key_0_683;
          put_stuckKeys_2_value_27 <= put_Key_1_687;
          put_stuckKeys_2_value_28 <= put_Key_2_691;
          put_stuckKeys_2_value_29 <= put_Key_3_695;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_735;
          put_stuckData_4_value_32 <= put_Data_0_686;
          put_stuckData_4_value_33 <= put_Data_1_690;
          put_stuckData_4_value_34 <= put_Data_2_694;
          put_stuckData_4_value_35 <= put_Data_3_698;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        434: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        435: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        436: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1755:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        437: begin
          put_stuckSize_6_index_37 <= put_childData_734;
          put_stuckSize_6_value_38 <= put_size_653;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childData_734;
          put_stuckKeys_2_value_26 <= put_Key_0_656;
          put_stuckKeys_2_value_27 <= put_Key_1_660;
          put_stuckKeys_2_value_28 <= put_Key_2_664;
          put_stuckKeys_2_value_29 <= put_Key_3_668;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childData_734;
          put_stuckData_4_value_32 <= put_Data_0_659;
          put_stuckData_4_value_33 <= put_Data_1_663;
          put_stuckData_4_value_34 <= put_Data_2_667;
          put_stuckData_4_value_35 <= put_Data_3_671;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1756:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        438: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1756:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        439: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1756:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        440: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1756:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        441: begin
          case (put_size_626)
            0: begin
              put_Key_0_629 <= put_midKey_737;
              put_Data_0_632 <= put_indexLeft_735;
            end
            1: begin
              put_Key_1_633 <= put_midKey_737;
              put_Data_1_636 <= put_indexLeft_735;
            end
            2: begin
              put_Key_2_637 <= put_midKey_737;
              put_Data_2_640 <= put_indexLeft_735;
            end
            3: begin
              put_Key_3_641 <= put_midKey_737;
              put_Data_3_644 <= put_indexLeft_735;
            end
          endcase
          put_size_626 <= put_size_626+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0423:<init>|  Btree.java:0422:Push|  Btree.java:1758:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        442: begin
          case (put_size_626)
            0: begin
              put_Key_0_629 <= put_midKey_737;
              put_Data_0_632 <= put_childData_734;
            end
            1: begin
              put_Key_1_633 <= put_midKey_737;
              put_Data_1_636 <= put_childData_734;
            end
            2: begin
              put_Key_2_637 <= put_midKey_737;
              put_Data_2_640 <= put_childData_734;
            end
            3: begin
              put_Key_3_641 <= put_midKey_737;
              put_Data_3_644 <= put_childData_734;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0480:<init>|  Btree.java:0479:SetPastLastElement|  Btree.java:1759:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        443: begin
          put_stuckSize_6_index_37 <= put_index_625;
          put_stuckSize_6_value_38 <= put_size_626;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_625;
          put_stuckKeys_2_value_26 <= put_Key_0_629;
          put_stuckKeys_2_value_27 <= put_Key_1_633;
          put_stuckKeys_2_value_28 <= put_Key_2_637;
          put_stuckKeys_2_value_29 <= put_Key_3_641;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_625;
          put_stuckData_4_value_32 <= put_Data_0_632;
          put_stuckData_4_value_33 <= put_Data_1_636;
          put_stuckData_4_value_34 <= put_Data_2_640;
          put_stuckData_4_value_35 <= put_Data_3_644;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1760:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        444: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1760:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        445: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1760:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        446: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1760:splitBranchAtTop|  Btree.java:2403:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Then|  Chip.java:0610:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        447: begin
          put_pc <= 449;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        448: begin
          put_parent_104 <= put_child_103;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2408:Else|  Chip.java:0620:<init>|  Btree.java:2397:<init>|  Btree.java:2396:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        449: begin
          put_pc <= 199;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2412:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2374:<init>|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2358:<init>|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2332:<init>|  Btree.java:2331:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        450: begin
          put_position_769 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2434:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        451: begin
          put_index_742 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        452: begin
          put_stuckSize_5_index_36 <= put_index_742;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_742;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_742;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_742;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        453: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        454: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        455: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        456: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        457: begin
          put_size_743 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_744 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_746 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_749 <= stuckData_stuckData_3_result_0;
          put_Key_1_750 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_753 <= stuckData_stuckData_3_result_1;
          put_Key_2_754 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_757 <= stuckData_stuckData_3_result_2;
          put_Key_3_758 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_761 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2436:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        458: begin
          if (put_isLeaf_744 == 0) begin
            put_pc <= 461;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2439:<init>|  Btree.java:2438:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        459: begin
          put_pc <= 982;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2440:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2439:<init>|  Btree.java:2438:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        460: begin
          put_pc <= 461;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2439:<init>|  Btree.java:2438:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        461: begin
          put_success_860 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1813:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        462: begin
          put_index_774 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        463: begin
          put_stuckSize_5_index_36 <= put_index_774;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_774;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_774;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_774;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        464: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        465: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        466: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        467: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        468: begin
          put_size_775 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_776 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_778 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_781 <= stuckData_stuckData_3_result_0;
          put_Key_1_782 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_785 <= stuckData_stuckData_3_result_1;
          put_Key_2_786 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_789 <= stuckData_stuckData_3_result_2;
          put_Key_3_790 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_793 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:1814:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        469: begin
          put_test_861 <= put_size_775==1 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0785:<init>|  Chip.java:0785:Eq|  Btree.java:1816:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        470: begin
          if (put_test_861 == 0) begin
            put_pc <= 522;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0585:<init>|  Chip.java:0584:GOZero|  Btree.java:1817:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        471: begin
          put_indexLeft_857 <= put_Data_0_781;
          put_indexRight_858 <= put_Data_1_785;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1820:<init>|  Btree.java:1819:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        472: begin
          put_index_801 <= put_indexLeft_857;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        473: begin
          put_stuckSize_5_index_36 <= put_index_801;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_801;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_801;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_801;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        474: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        475: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        476: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        477: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        478: begin
          put_size_802 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_803 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_805 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_808 <= stuckData_stuckData_3_result_0;
          put_Key_1_809 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_812 <= stuckData_stuckData_3_result_1;
          put_Key_2_813 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_816 <= stuckData_stuckData_3_result_2;
          put_Key_3_817 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_820 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1830:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        479: begin
          put_index_828 <= put_indexRight_858;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        480: begin
          put_stuckSize_5_index_36 <= put_index_828;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_828;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_828;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_828;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        481: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        482: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        483: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        484: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        485: begin
          put_size_829 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_830 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_832 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_835 <= stuckData_stuckData_3_result_0;
          put_Key_1_836 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_839 <= stuckData_stuckData_3_result_1;
          put_Key_2_840 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_843 <= stuckData_stuckData_3_result_2;
          put_Key_3_844 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_847 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1831:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        486: begin
          if (put_isLeaf_803 == 0) begin
            put_pc <= 522;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        487: begin
          if (put_isLeaf_830 == 0) begin
            put_pc <= 521;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        488: begin
          put_MergeSuccess_800 <= 0;
          case (put_size_802)
            0: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                4: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1251:<init>|  Btree.java:1250:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        489: begin
          if (put_MergeSuccess_800 == 0) begin
            put_pc <= 493;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        490: begin
          put_MergeSuccess_800 <= 0;
          case (put_size_775)
            0: begin
              case (put_size_802)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_0_778 <= put_Key_0_805;
                  put_Data_0_781 <= put_Data_0_808;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_Key_0_778 <= put_Key_0_805;
                  put_Data_0_781 <= put_Data_0_808;
                  put_Key_1_782 <= put_Key_1_809;
                  put_Data_1_785 <= put_Data_1_812;
                  put_size_775 <= put_size_775 + 2;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                  put_Key_0_778 <= put_Key_0_805;
                  put_Data_0_781 <= put_Data_0_808;
                  put_Key_1_782 <= put_Key_1_809;
                  put_Data_1_785 <= put_Data_1_812;
                  put_Key_2_786 <= put_Key_2_813;
                  put_Data_2_789 <= put_Data_2_816;
                  put_size_775 <= put_size_775 + 3;
                  put_MergeSuccess_800 <= 1;
                end
                4: begin
                  put_Key_0_778 <= put_Key_0_805;
                  put_Data_0_781 <= put_Data_0_808;
                  put_Key_1_782 <= put_Key_1_809;
                  put_Data_1_785 <= put_Data_1_812;
                  put_Key_2_786 <= put_Key_2_813;
                  put_Data_2_789 <= put_Data_2_816;
                  put_Key_3_790 <= put_Key_3_817;
                  put_Data_3_793 <= put_Data_3_820;
                  put_size_775 <= put_size_775 + 4;
                  put_MergeSuccess_800 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_802)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_1_782 <= put_Key_0_805;
                  put_Data_1_785 <= put_Data_0_808;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_Key_1_782 <= put_Key_0_805;
                  put_Data_1_785 <= put_Data_0_808;
                  put_Key_2_786 <= put_Key_1_809;
                  put_Data_2_789 <= put_Data_1_812;
                  put_size_775 <= put_size_775 + 2;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                  put_Key_1_782 <= put_Key_0_805;
                  put_Data_1_785 <= put_Data_0_808;
                  put_Key_2_786 <= put_Key_1_809;
                  put_Data_2_789 <= put_Data_1_812;
                  put_Key_3_790 <= put_Key_2_813;
                  put_Data_3_793 <= put_Data_2_816;
                  put_size_775 <= put_size_775 + 3;
                  put_MergeSuccess_800 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_802)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_2_786 <= put_Key_0_805;
                  put_Data_2_789 <= put_Data_0_808;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_Key_2_786 <= put_Key_0_805;
                  put_Data_2_789 <= put_Data_0_808;
                  put_Key_3_790 <= put_Key_1_809;
                  put_Data_3_793 <= put_Data_1_812;
                  put_size_775 <= put_size_775 + 2;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_802)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_3_790 <= put_Key_0_805;
                  put_Data_3_793 <= put_Data_0_808;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_802)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1279:Then|  Chip.java:0610:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        491: begin
          put_MergeSuccess_800 <= 0;
          case (put_size_775)
            0: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_0_778 <= put_Key_0_832;
                  put_Data_0_781 <= put_Data_0_835;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_Key_0_778 <= put_Key_0_832;
                  put_Data_0_781 <= put_Data_0_835;
                  put_Key_1_782 <= put_Key_1_836;
                  put_Data_1_785 <= put_Data_1_839;
                  put_size_775 <= put_size_775 + 2;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                  put_Key_0_778 <= put_Key_0_832;
                  put_Data_0_781 <= put_Data_0_835;
                  put_Key_1_782 <= put_Key_1_836;
                  put_Data_1_785 <= put_Data_1_839;
                  put_Key_2_786 <= put_Key_2_840;
                  put_Data_2_789 <= put_Data_2_843;
                  put_size_775 <= put_size_775 + 3;
                  put_MergeSuccess_800 <= 1;
                end
                4: begin
                  put_Key_0_778 <= put_Key_0_832;
                  put_Data_0_781 <= put_Data_0_835;
                  put_Key_1_782 <= put_Key_1_836;
                  put_Data_1_785 <= put_Data_1_839;
                  put_Key_2_786 <= put_Key_2_840;
                  put_Data_2_789 <= put_Data_2_843;
                  put_Key_3_790 <= put_Key_3_844;
                  put_Data_3_793 <= put_Data_3_847;
                  put_size_775 <= put_size_775 + 4;
                  put_MergeSuccess_800 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_1_782 <= put_Key_0_832;
                  put_Data_1_785 <= put_Data_0_835;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_Key_1_782 <= put_Key_0_832;
                  put_Data_1_785 <= put_Data_0_835;
                  put_Key_2_786 <= put_Key_1_836;
                  put_Data_2_789 <= put_Data_1_839;
                  put_size_775 <= put_size_775 + 2;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                  put_Key_1_782 <= put_Key_0_832;
                  put_Data_1_785 <= put_Data_0_835;
                  put_Key_2_786 <= put_Key_1_836;
                  put_Data_2_789 <= put_Data_1_839;
                  put_Key_3_790 <= put_Key_2_840;
                  put_Data_3_793 <= put_Data_2_843;
                  put_size_775 <= put_size_775 + 3;
                  put_MergeSuccess_800 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_2_786 <= put_Key_0_832;
                  put_Data_2_789 <= put_Data_0_835;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                  put_Key_2_786 <= put_Key_0_832;
                  put_Data_2_789 <= put_Data_0_835;
                  put_Key_3_790 <= put_Key_1_836;
                  put_Data_3_793 <= put_Data_1_839;
                  put_size_775 <= put_size_775 + 2;
                  put_MergeSuccess_800 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                  put_Key_3_790 <= put_Key_0_832;
                  put_Data_3_793 <= put_Data_0_835;
                  put_size_775 <= put_size_775 + 1;
                  put_MergeSuccess_800 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_829)
                0: begin
                  put_size_775 <= put_size_775 + 0;
                  put_MergeSuccess_800 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1280:Then|  Chip.java:0610:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        492: begin
          put_pc <= 493;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1278:<init>|  Btree.java:1277:merge|  Btree.java:1837:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        493: begin
          if (put_MergeSuccess_800 == 0) begin
            put_pc <= 520;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        494: begin
          put_isLeaf_776 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1840:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        495: begin
          put_stuckSize_6_index_37 <= put_index_774;
          put_stuckSize_6_value_38 <= put_size_775;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_index_774;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_776;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_774;
          put_stuckKeys_2_value_26 <= put_Key_0_778;
          put_stuckKeys_2_value_27 <= put_Key_1_782;
          put_stuckKeys_2_value_28 <= put_Key_2_786;
          put_stuckKeys_2_value_29 <= put_Key_3_790;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_774;
          put_stuckData_4_value_32 <= put_Data_0_781;
          put_stuckData_4_value_33 <= put_Data_1_785;
          put_stuckData_4_value_34 <= put_Data_2_789;
          put_stuckData_4_value_35 <= put_Data_3_793;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        496: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        497: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        498: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        499: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1841:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        500: begin
          put_root_863 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        501: begin
          put_freeNext_9_index_194 <= put_root_863;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        502: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        503: begin
          put_next_862 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_863;
          put_freeNext_10_value_196 <= put_indexLeft_857;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_864 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        504: begin
          put_stuckIsFree_11_index_197 <= put_indexLeft_857;
          put_stuckIsFree_11_value_198 <= put_isFree_864;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        505: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        506: begin
          put_freeNext_10_index_195 <= put_indexLeft_857;
          put_freeNext_10_value_196 <= put_next_862;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        507: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        508: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        509: begin
          put_root_866 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        510: begin
          put_freeNext_9_index_194 <= put_root_866;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        511: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        512: begin
          put_next_865 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_866;
          put_freeNext_10_value_196 <= put_indexRight_858;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_867 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        513: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_858;
          put_stuckIsFree_11_value_198 <= put_isFree_867;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        514: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        515: begin
          put_freeNext_10_index_195 <= put_indexRight_858;
          put_freeNext_10_value_196 <= put_next_865;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        516: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        517: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1842:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        518: begin
          put_success_860 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1843:Then|  Chip.java:0610:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        519: begin
          put_pc <= 520;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1839:<init>|  Btree.java:1838:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        520: begin
          put_pc <= 521;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1836:<init>|  Btree.java:1835:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        521: begin
          put_pc <= 522;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1834:<init>|  Btree.java:1833:code|  Chip.java:0530:<init>|  Btree.java:1812:<init>|  Btree.java:1811:mergeLeavesIntoRoot|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        522: begin
          if (put_success_860 == 0) begin
            put_pc <= 525;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2444:<init>|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        523: begin
          put_pc <= 982;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2445:Then|  Chip.java:0610:<init>|  Btree.java:2444:<init>|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        524: begin
          put_pc <= 525;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2444:<init>|  Btree.java:2443:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        525: begin
          put_index_868 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        526: begin
          put_stuckSize_5_index_36 <= put_index_868;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_868;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_868;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_868;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        527: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        528: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        529: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        530: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        531: begin
          put_size_869 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_870 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_872 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_875 <= stuckData_stuckData_3_result_0;
          put_Key_1_876 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_879 <= stuckData_stuckData_3_result_1;
          put_Key_2_880 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_883 <= stuckData_stuckData_3_result_2;
          put_Key_3_884 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_887 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2018:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        532: begin
          put_success_956 <= 0;
          if (put_size_869 != 1) begin
            put_pc <= 578;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:2023:<init>|  Btree.java:2022:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        533: begin
          put_midKey_955 <= put_Key_0_872;
          put_indexLeft_953 <= put_Data_0_875;
          put_indexRight_954 <= put_Data_1_879;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2041:<init>|  Btree.java:2040:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        534: begin
          if (put_isLeaf_897 == 0) begin
            put_pc <= 536;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        535: begin
          put_pc <= 578;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        536: begin
          if (put_isLeaf_924 == 0) begin
            put_pc <= 538;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        537: begin
          put_pc <= 578;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        538: begin
          put_index_895 <= put_indexLeft_953;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        539: begin
          put_stuckSize_5_index_36 <= put_index_895;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_895;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_895;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_895;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        540: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        541: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        542: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        543: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        544: begin
          put_size_896 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_897 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_899 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_902 <= stuckData_stuckData_3_result_0;
          put_Key_1_903 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_906 <= stuckData_stuckData_3_result_1;
          put_Key_2_907 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_910 <= stuckData_stuckData_3_result_2;
          put_Key_3_911 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_914 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2057:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        545: begin
          put_index_922 <= put_indexRight_954;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        546: begin
          put_stuckSize_5_index_36 <= put_index_922;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_922;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_922;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_922;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        547: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        548: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        549: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        550: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        551: begin
          put_size_923 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_924 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_926 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_929 <= stuckData_stuckData_3_result_0;
          put_Key_1_930 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_933 <= stuckData_stuckData_3_result_1;
          put_Key_2_934 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_937 <= stuckData_stuckData_3_result_2;
          put_Key_3_938 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_941 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2058:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        552: begin
          put_MergeSuccess_894 <= 0;
          case (put_size_896)
            0: begin
              case (put_size_923)
                0: begin
                  put_Key_0_872 <= put_midKey_955;
                  put_Data_0_875 <= put_Data_0_902;
                  put_Data_1_879 <= put_Data_0_929;
                  put_size_869 <= 1;
                  put_MergeSuccess_894 <= 1;
                end
                1: begin
                  put_Key_0_872 <= put_midKey_955;
                  put_Data_0_875 <= put_Data_0_902;
                  put_Key_1_876 <= put_Key_0_926;
                  put_Data_1_879 <= put_Data_0_929;
                  put_Data_2_883 <= put_Data_1_933;
                  put_size_869 <= 2;
                  put_MergeSuccess_894 <= 1;
                end
                2: begin
                  put_Key_0_872 <= put_midKey_955;
                  put_Data_0_875 <= put_Data_0_902;
                  put_Key_1_876 <= put_Key_0_926;
                  put_Data_1_879 <= put_Data_0_929;
                  put_Key_2_880 <= put_Key_1_930;
                  put_Data_2_883 <= put_Data_1_933;
                  put_Data_3_887 <= put_Data_2_937;
                  put_size_869 <= 3;
                  put_MergeSuccess_894 <= 1;
                end
                3: begin
                end
              endcase
            end
            1: begin
              case (put_size_923)
                0: begin
                  put_Key_0_872 <= put_Key_0_899;
                  put_Data_0_875 <= put_Data_0_902;
                  put_Key_1_876 <= put_midKey_955;
                  put_Data_1_879 <= put_Data_1_906;
                  put_Data_2_883 <= put_Data_0_929;
                  put_size_869 <= 2;
                  put_MergeSuccess_894 <= 1;
                end
                1: begin
                  put_Key_0_872 <= put_Key_0_899;
                  put_Data_0_875 <= put_Data_0_902;
                  put_Key_1_876 <= put_midKey_955;
                  put_Data_1_879 <= put_Data_1_906;
                  put_Key_2_880 <= put_Key_0_926;
                  put_Data_2_883 <= put_Data_0_929;
                  put_Data_3_887 <= put_Data_1_933;
                  put_size_869 <= 3;
                  put_MergeSuccess_894 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (put_size_923)
                0: begin
                  put_Key_0_872 <= put_Key_0_899;
                  put_Data_0_875 <= put_Data_0_902;
                  put_Key_1_876 <= put_Key_1_903;
                  put_Data_1_879 <= put_Data_1_906;
                  put_Key_2_880 <= put_midKey_955;
                  put_Data_2_883 <= put_Data_2_910;
                  put_Data_3_887 <= put_Data_0_929;
                  put_size_869 <= 3;
                  put_MergeSuccess_894 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            3: begin
              case (put_size_923)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1329:<init>|  Btree.java:1328:mergeButOne|  Btree.java:2059:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        553: begin
          if (put_MergeSuccess_894 == 0) begin
            put_pc <= 578;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        554: begin
          put_stuckSize_6_index_37 <= put_index_868;
          put_stuckSize_6_value_38 <= put_size_869;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_868;
          put_stuckKeys_2_value_26 <= put_Key_0_872;
          put_stuckKeys_2_value_27 <= put_Key_1_876;
          put_stuckKeys_2_value_28 <= put_Key_2_880;
          put_stuckKeys_2_value_29 <= put_Key_3_884;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_868;
          put_stuckData_4_value_32 <= put_Data_0_875;
          put_stuckData_4_value_33 <= put_Data_1_879;
          put_stuckData_4_value_34 <= put_Data_2_883;
          put_stuckData_4_value_35 <= put_Data_3_887;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        555: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        556: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        557: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2062:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        558: begin
          put_root_959 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        559: begin
          put_freeNext_9_index_194 <= put_root_959;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        560: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        561: begin
          put_next_958 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_959;
          put_freeNext_10_value_196 <= put_indexLeft_953;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_960 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        562: begin
          put_stuckIsFree_11_index_197 <= put_indexLeft_953;
          put_stuckIsFree_11_value_198 <= put_isFree_960;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        563: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        564: begin
          put_freeNext_10_index_195 <= put_indexLeft_953;
          put_freeNext_10_value_196 <= put_next_958;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        565: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        566: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        567: begin
          put_root_962 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        568: begin
          put_freeNext_9_index_194 <= put_root_962;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        569: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        570: begin
          put_next_961 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_962;
          put_freeNext_10_value_196 <= put_indexRight_954;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_963 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        571: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_954;
          put_stuckIsFree_11_value_198 <= put_isFree_963;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        572: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        573: begin
          put_freeNext_10_index_195 <= put_indexRight_954;
          put_freeNext_10_value_196 <= put_next_961;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        574: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        575: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2063:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        576: begin
          put_success_956 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2064:Then|  Chip.java:0610:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        577: begin
          put_pc <= 578;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2061:<init>|  Btree.java:2060:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2056:<init>|  Btree.java:2055:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2054:<init>|  Btree.java:2053:code|  Chip.java:0530:<init>|  Btree.java:2021:<init>|  Btree.java:2020:mergeBranchesIntoRoot|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        578: begin
          if (put_success_956 == 0) begin
            put_pc <= 587;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        579: begin
          put_index_742 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0266:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        580: begin
          put_stuckSize_5_index_36 <= put_index_742;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_742;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_742;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_742;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        581: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        582: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        583: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        584: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        585: begin
          put_size_743 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_744 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_746 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_749 <= stuckData_stuckData_3_result_0;
          put_Key_1_750 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_753 <= stuckData_stuckData_3_result_1;
          put_Key_2_754 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_757 <= stuckData_stuckData_3_result_2;
          put_Key_3_758 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_761 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0267:stuckGetRoot|  Btree.java:2451:Then|  Chip.java:0610:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        586: begin
          put_pc <= 587;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2450:<init>|  Btree.java:2449:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        587: begin
          put_success_1024 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1941:<init>|  Btree.java:1940:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        588: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 630;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1949:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        589: begin
          put_size_1019 <= put_size_743;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1950:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        590: begin
          case (put_size_1019)
            1: begin
              put_indexLeft_1021 <= put_Data_0_749;
              put_indexRight_1022 <= put_Data_1_753;
            end
            2: begin
              put_indexLeft_1021 <= put_Data_1_753;
              put_indexRight_1022 <= put_Data_2_757;
            end
            3: begin
              put_indexLeft_1021 <= put_Data_2_757;
              put_indexRight_1022 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1953:<init>|  Btree.java:1952:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        591: begin
          put_index_964 <= put_indexLeft_1021;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        592: begin
          put_stuckSize_5_index_36 <= put_index_964;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_964;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_964;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_964;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        593: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        594: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        595: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        596: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        597: begin
          put_size_965 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_966 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_968 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_971 <= stuckData_stuckData_3_result_0;
          put_Key_1_972 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_975 <= stuckData_stuckData_3_result_1;
          put_Key_2_976 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_979 <= stuckData_stuckData_3_result_2;
          put_Key_3_980 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_983 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1967:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        598: begin
          put_index_991 <= put_indexRight_1022;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        599: begin
          put_stuckSize_5_index_36 <= put_index_991;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_991;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_991;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_991;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        600: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        601: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        602: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        603: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        604: begin
          put_size_992 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_993 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_995 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_998 <= stuckData_stuckData_3_result_0;
          put_Key_1_999 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1002 <= stuckData_stuckData_3_result_1;
          put_Key_2_1003 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1006 <= stuckData_stuckData_3_result_2;
          put_Key_3_1007 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1010 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1968:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        605: begin
          if (put_isLeaf_966 == 0) begin
            put_pc <= 630;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        606: begin
          if (put_isLeaf_993 == 0) begin
            put_pc <= 629;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        607: begin
          put_MergeSuccess_990 <= 0;
          case (put_size_965)
            0: begin
              case (put_size_992)
                0: begin
                  put_size_965 <= put_size_965 + 0;
                  put_MergeSuccess_990 <= 1;
                end
                1: begin
                  put_Key_0_968 <= put_Key_0_995;
                  put_Data_0_971 <= put_Data_0_998;
                  put_size_965 <= put_size_965 + 1;
                  put_MergeSuccess_990 <= 1;
                end
                2: begin
                  put_Key_0_968 <= put_Key_0_995;
                  put_Data_0_971 <= put_Data_0_998;
                  put_Key_1_972 <= put_Key_1_999;
                  put_Data_1_975 <= put_Data_1_1002;
                  put_size_965 <= put_size_965 + 2;
                  put_MergeSuccess_990 <= 1;
                end
                3: begin
                  put_Key_0_968 <= put_Key_0_995;
                  put_Data_0_971 <= put_Data_0_998;
                  put_Key_1_972 <= put_Key_1_999;
                  put_Data_1_975 <= put_Data_1_1002;
                  put_Key_2_976 <= put_Key_2_1003;
                  put_Data_2_979 <= put_Data_2_1006;
                  put_size_965 <= put_size_965 + 3;
                  put_MergeSuccess_990 <= 1;
                end
                4: begin
                  put_Key_0_968 <= put_Key_0_995;
                  put_Data_0_971 <= put_Data_0_998;
                  put_Key_1_972 <= put_Key_1_999;
                  put_Data_1_975 <= put_Data_1_1002;
                  put_Key_2_976 <= put_Key_2_1003;
                  put_Data_2_979 <= put_Data_2_1006;
                  put_Key_3_980 <= put_Key_3_1007;
                  put_Data_3_983 <= put_Data_3_1010;
                  put_size_965 <= put_size_965 + 4;
                  put_MergeSuccess_990 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_992)
                0: begin
                  put_size_965 <= put_size_965 + 0;
                  put_MergeSuccess_990 <= 1;
                end
                1: begin
                  put_Key_1_972 <= put_Key_0_995;
                  put_Data_1_975 <= put_Data_0_998;
                  put_size_965 <= put_size_965 + 1;
                  put_MergeSuccess_990 <= 1;
                end
                2: begin
                  put_Key_1_972 <= put_Key_0_995;
                  put_Data_1_975 <= put_Data_0_998;
                  put_Key_2_976 <= put_Key_1_999;
                  put_Data_2_979 <= put_Data_1_1002;
                  put_size_965 <= put_size_965 + 2;
                  put_MergeSuccess_990 <= 1;
                end
                3: begin
                  put_Key_1_972 <= put_Key_0_995;
                  put_Data_1_975 <= put_Data_0_998;
                  put_Key_2_976 <= put_Key_1_999;
                  put_Data_2_979 <= put_Data_1_1002;
                  put_Key_3_980 <= put_Key_2_1003;
                  put_Data_3_983 <= put_Data_2_1006;
                  put_size_965 <= put_size_965 + 3;
                  put_MergeSuccess_990 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_992)
                0: begin
                  put_size_965 <= put_size_965 + 0;
                  put_MergeSuccess_990 <= 1;
                end
                1: begin
                  put_Key_2_976 <= put_Key_0_995;
                  put_Data_2_979 <= put_Data_0_998;
                  put_size_965 <= put_size_965 + 1;
                  put_MergeSuccess_990 <= 1;
                end
                2: begin
                  put_Key_2_976 <= put_Key_0_995;
                  put_Data_2_979 <= put_Data_0_998;
                  put_Key_3_980 <= put_Key_1_999;
                  put_Data_3_983 <= put_Data_1_1002;
                  put_size_965 <= put_size_965 + 2;
                  put_MergeSuccess_990 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_992)
                0: begin
                  put_size_965 <= put_size_965 + 0;
                  put_MergeSuccess_990 <= 1;
                end
                1: begin
                  put_Key_3_980 <= put_Key_0_995;
                  put_Data_3_983 <= put_Data_0_998;
                  put_size_965 <= put_size_965 + 1;
                  put_MergeSuccess_990 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_992)
                0: begin
                  put_size_965 <= put_size_965 + 0;
                  put_MergeSuccess_990 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1974:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        608: begin
          if (put_MergeSuccess_990 == 0) begin
            put_pc <= 628;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        609: begin
          put_size_743 <= put_size_743-1;
          put_success_1024 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1978:<init>|  Btree.java:1977:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        610: begin
          put_stuckSize_6_index_37 <= put_index_964;
          put_stuckSize_6_value_38 <= put_size_965;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_964;
          put_stuckKeys_2_value_26 <= put_Key_0_968;
          put_stuckKeys_2_value_27 <= put_Key_1_972;
          put_stuckKeys_2_value_28 <= put_Key_2_976;
          put_stuckKeys_2_value_29 <= put_Key_3_980;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_964;
          put_stuckData_4_value_32 <= put_Data_0_971;
          put_stuckData_4_value_33 <= put_Data_1_975;
          put_stuckData_4_value_34 <= put_Data_2_979;
          put_stuckData_4_value_35 <= put_Data_3_983;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        611: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        612: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        613: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1987:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        614: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        615: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        616: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        617: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1988:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        618: begin
          put_root_1027 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        619: begin
          put_freeNext_9_index_194 <= put_root_1027;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        620: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        621: begin
          put_next_1026 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1027;
          put_freeNext_10_value_196 <= put_indexRight_1022;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1028 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        622: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1022;
          put_stuckIsFree_11_value_198 <= put_isFree_1028;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        623: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        624: begin
          put_freeNext_10_index_195 <= put_indexRight_1022;
          put_freeNext_10_value_196 <= put_next_1026;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        625: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        626: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1989:Then|  Chip.java:0610:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        627: begin
          put_pc <= 628;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1976:<init>|  Btree.java:1975:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        628: begin
          put_pc <= 629;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1973:<init>|  Btree.java:1972:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        629: begin
          put_pc <= 630;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1971:<init>|  Btree.java:1970:code|  Chip.java:0530:<init>|  Btree.java:1948:<init>|  Btree.java:1947:mergeLeavesAtTop|  Btree.java:2457:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        630: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 675;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2183:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        631: begin
          put_success_1089 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2184:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        632: begin
          put_size_1084 <= put_size_743;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2185:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        633: begin
          case (put_size_1084)
            1: begin
              put_indexLeft_1086 <= put_Data_0_749;
              put_indexRight_1087 <= put_Data_1_753;
            end
            2: begin
              put_indexLeft_1086 <= put_Data_1_753;
              put_indexRight_1087 <= put_Data_2_757;
            end
            3: begin
              put_indexLeft_1086 <= put_Data_2_757;
              put_indexRight_1087 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2188:<init>|  Btree.java:2187:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        634: begin
          put_index_1029 <= put_indexLeft_1086;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        635: begin
          put_stuckSize_5_index_36 <= put_index_1029;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1029;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1029;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1029;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        636: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        637: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        638: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        639: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        640: begin
          put_size_1030 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1031 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1033 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1036 <= stuckData_stuckData_3_result_0;
          put_Key_1_1037 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1040 <= stuckData_stuckData_3_result_1;
          put_Key_2_1041 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1044 <= stuckData_stuckData_3_result_2;
          put_Key_3_1045 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1048 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        641: begin
          put_index_1056 <= put_indexRight_1087;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        642: begin
          put_stuckSize_5_index_36 <= put_index_1056;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1056;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1056;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1056;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        643: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        644: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        645: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        646: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        647: begin
          put_size_1057 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1058 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1060 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1063 <= stuckData_stuckData_3_result_0;
          put_Key_1_1064 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1067 <= stuckData_stuckData_3_result_1;
          put_Key_2_1068 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1071 <= stuckData_stuckData_3_result_2;
          put_Key_3_1072 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1075 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        648: begin
          if (put_isLeaf_1031 == 0) begin
            put_pc <= 650;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        649: begin
          put_pc <= 675;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        650: begin
          if (put_isLeaf_1058 == 0) begin
            put_pc <= 652;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        651: begin
          put_pc <= 675;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        652: begin
          case (put_size_743)
            1: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            2: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            3: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            4: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_size_743 <= put_size_743-1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0452:<init>|  Btree.java:0451:Pop|  Btree.java:2209:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        653: begin
          put_MergeSuccess_1055 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2210:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        654: begin
          case (put_size_1030)
            0: begin
              case (put_size_1057)
                0: begin
                  put_Key_0_1033 <= put_Key_763;
                  put_Data_1_1040 <= put_Data_0_1063;
                  put_size_1030 <= put_size_1030 + 1;
                  put_MergeSuccess_1055 <= 1;
                end
                1: begin
                  put_Key_0_1033 <= put_Key_763;
                  put_Key_1_1037 <= put_Key_0_1060;
                  put_Data_1_1040 <= put_Data_0_1063;
                  put_Data_2_1044 <= put_Data_1_1067;
                  put_size_1030 <= put_size_1030 + 2;
                  put_MergeSuccess_1055 <= 1;
                end
                2: begin
                  put_Key_0_1033 <= put_Key_763;
                  put_Key_1_1037 <= put_Key_0_1060;
                  put_Data_1_1040 <= put_Data_0_1063;
                  put_Key_2_1041 <= put_Key_1_1064;
                  put_Data_2_1044 <= put_Data_1_1067;
                  put_Data_3_1048 <= put_Data_2_1071;
                  put_size_1030 <= put_size_1030 + 3;
                  put_MergeSuccess_1055 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (put_size_1057)
                0: begin
                  put_Key_1_1037 <= put_Key_763;
                  put_Data_2_1044 <= put_Data_0_1063;
                  put_size_1030 <= put_size_1030 + 1;
                  put_MergeSuccess_1055 <= 1;
                end
                1: begin
                  put_Key_1_1037 <= put_Key_763;
                  put_Key_2_1041 <= put_Key_0_1060;
                  put_Data_2_1044 <= put_Data_0_1063;
                  put_Data_3_1048 <= put_Data_1_1067;
                  put_size_1030 <= put_size_1030 + 2;
                  put_MergeSuccess_1055 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1057)
                0: begin
                  put_Key_2_1041 <= put_Key_763;
                  put_Data_3_1048 <= put_Data_0_1063;
                  put_size_1030 <= put_size_1030 + 1;
                  put_MergeSuccess_1055 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1057)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1057)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2210:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        655: begin
          if (put_MergeSuccess_1055 == 0) begin
            put_pc <= 675;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        656: begin
          put_success_1089 <= 1;
          case (put_size_743)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1086;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1086;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1086;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1086;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2214:<init>|  Btree.java:2213:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        657: begin
          put_stuckSize_6_index_37 <= put_index_1029;
          put_stuckSize_6_value_38 <= put_size_1030;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1029;
          put_stuckKeys_2_value_26 <= put_Key_0_1033;
          put_stuckKeys_2_value_27 <= put_Key_1_1037;
          put_stuckKeys_2_value_28 <= put_Key_2_1041;
          put_stuckKeys_2_value_29 <= put_Key_3_1045;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1029;
          put_stuckData_4_value_32 <= put_Data_0_1036;
          put_stuckData_4_value_33 <= put_Data_1_1040;
          put_stuckData_4_value_34 <= put_Data_2_1044;
          put_stuckData_4_value_35 <= put_Data_3_1048;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        658: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        659: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        660: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        661: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        662: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        663: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        664: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        665: begin
          put_root_1092 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        666: begin
          put_freeNext_9_index_194 <= put_root_1092;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        667: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        668: begin
          put_next_1091 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1092;
          put_freeNext_10_value_196 <= put_indexRight_1087;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1093 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        669: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1087;
          put_stuckIsFree_11_value_198 <= put_isFree_1093;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        670: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        671: begin
          put_freeNext_10_index_195 <= put_indexRight_1087;
          put_freeNext_10_value_196 <= put_next_1091;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        672: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        673: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        674: begin
          put_pc <= 675;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:2458:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        675: begin
          put_KeyCompares_0_747 <= put_k_0 <= put_Key_0_746 && 0 < put_size_743;
          put_KeyCollapse_0_748 <= 0;
          put_KeyCompares_1_751 <= put_k_0 >  put_Key_0_746 && put_k_0 <= put_Key_1_750 && 1 < put_size_743;
          put_KeyCollapse_1_752 <= 1;
          put_KeyCompares_2_755 <= put_k_0 >  put_Key_1_750 && put_k_0 <= put_Key_2_754 && 2 < put_size_743;
          put_KeyCollapse_2_756 <= 2;
          put_KeyCompares_3_759 <= put_k_0 >  put_Key_2_754 && put_k_0 <= put_Key_3_758 && 3 < put_size_743;
          put_KeyCollapse_3_760 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        676: begin
          if (put_KeyCompares_1_751) begin
            put_KeyCompares_0_747 <= 1;
            put_KeyCollapse_0_748 <= put_KeyCollapse_1_752;
          end
          if (put_KeyCompares_3_759) begin
            put_KeyCompares_2_755 <= 1;
            put_KeyCollapse_2_756 <= put_KeyCollapse_3_760;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        677: begin
          if (put_KeyCompares_2_755) begin
            put_KeyCompares_0_747 <= 1;
            put_KeyCollapse_0_748 <= put_KeyCollapse_2_756;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        678: begin
          if (put_KeyCompares_0_747) begin
            put_Found_762 <= 1;
            case (put_KeyCollapse_0_748)
              0: begin
                put_StuckIndex_767 <= 0;
                put_FoundKey_764 <= put_Key_0_746;
                put_Data_765 <= put_Data_0_749;
              end
              1: begin
                put_StuckIndex_767 <= 1;
                put_FoundKey_764 <= put_Key_1_750;
                put_Data_765 <= put_Data_1_753;
              end
              2: begin
                put_StuckIndex_767 <= 2;
                put_FoundKey_764 <= put_Key_2_754;
                put_Data_765 <= put_Data_2_757;
              end
              3: begin
                put_StuckIndex_767 <= 3;
                put_FoundKey_764 <= put_Key_3_758;
                put_Data_765 <= put_Data_3_761;
              end
            endcase
          end
          else begin
            put_Found_762 <= 0;
            case (put_size_743)
              0: begin
                put_StuckIndex_767 <= 0;
                put_Data_765 <= put_Data_0_749;
              end
              1: begin
                put_StuckIndex_767 <= 1;
                put_Data_765 <= put_Data_1_753;
              end
              2: begin
                put_StuckIndex_767 <= 2;
                put_Data_765 <= put_Data_2_757;
              end
              3: begin
                put_StuckIndex_767 <= 3;
                put_Data_765 <= put_Data_3_761;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2459:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        679: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2461:<init>|  Btree.java:2460:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        680: begin
          if (put_Found_762 == 0) begin
            put_pc <= 959;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        681: begin
          if (put_StuckIndex_767 == 0) begin
            put_pc <= 867;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        682: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 726;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        683: begin
          case (put_StuckIndex_767)
            0: begin
              put_indexLeft_1150 <= put_Data_0_749;
              put_indexRight_1151 <= put_Data_1_753;
            end
            1: begin
              put_indexLeft_1150 <= put_Data_1_753;
              put_indexRight_1151 <= put_Data_2_757;
            end
            2: begin
              put_indexLeft_1150 <= put_Data_2_757;
              put_indexRight_1151 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        684: begin
          put_index_1094 <= put_indexLeft_1150;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        685: begin
          put_stuckSize_5_index_36 <= put_index_1094;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1094;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1094;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1094;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        686: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        687: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        688: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        689: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        690: begin
          put_size_1095 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1096 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1098 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1101 <= stuckData_stuckData_3_result_0;
          put_Key_1_1102 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1105 <= stuckData_stuckData_3_result_1;
          put_Key_2_1106 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1109 <= stuckData_stuckData_3_result_2;
          put_Key_3_1110 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1113 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        691: begin
          put_index_1121 <= put_indexRight_1151;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        692: begin
          put_stuckSize_5_index_36 <= put_index_1121;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1121;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1121;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1121;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        693: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        694: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        695: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        696: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        697: begin
          put_size_1122 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1123 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1125 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1128 <= stuckData_stuckData_3_result_0;
          put_Key_1_1129 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1132 <= stuckData_stuckData_3_result_1;
          put_Key_2_1133 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1136 <= stuckData_stuckData_3_result_2;
          put_Key_3_1137 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1140 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        698: begin
          if (put_isLeaf_1096 == 0) begin
            put_pc <= 726;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        699: begin
          if (put_isLeaf_1123 == 0) begin
            put_pc <= 725;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        700: begin
          put_MergeSuccess_1120 <= 0;
          case (put_size_1095)
            0: begin
              case (put_size_1122)
                0: begin
                  put_size_1095 <= put_size_1095 + 0;
                  put_MergeSuccess_1120 <= 1;
                end
                1: begin
                  put_Key_0_1098 <= put_Key_0_1125;
                  put_Data_0_1101 <= put_Data_0_1128;
                  put_size_1095 <= put_size_1095 + 1;
                  put_MergeSuccess_1120 <= 1;
                end
                2: begin
                  put_Key_0_1098 <= put_Key_0_1125;
                  put_Data_0_1101 <= put_Data_0_1128;
                  put_Key_1_1102 <= put_Key_1_1129;
                  put_Data_1_1105 <= put_Data_1_1132;
                  put_size_1095 <= put_size_1095 + 2;
                  put_MergeSuccess_1120 <= 1;
                end
                3: begin
                  put_Key_0_1098 <= put_Key_0_1125;
                  put_Data_0_1101 <= put_Data_0_1128;
                  put_Key_1_1102 <= put_Key_1_1129;
                  put_Data_1_1105 <= put_Data_1_1132;
                  put_Key_2_1106 <= put_Key_2_1133;
                  put_Data_2_1109 <= put_Data_2_1136;
                  put_size_1095 <= put_size_1095 + 3;
                  put_MergeSuccess_1120 <= 1;
                end
                4: begin
                  put_Key_0_1098 <= put_Key_0_1125;
                  put_Data_0_1101 <= put_Data_0_1128;
                  put_Key_1_1102 <= put_Key_1_1129;
                  put_Data_1_1105 <= put_Data_1_1132;
                  put_Key_2_1106 <= put_Key_2_1133;
                  put_Data_2_1109 <= put_Data_2_1136;
                  put_Key_3_1110 <= put_Key_3_1137;
                  put_Data_3_1113 <= put_Data_3_1140;
                  put_size_1095 <= put_size_1095 + 4;
                  put_MergeSuccess_1120 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_1122)
                0: begin
                  put_size_1095 <= put_size_1095 + 0;
                  put_MergeSuccess_1120 <= 1;
                end
                1: begin
                  put_Key_1_1102 <= put_Key_0_1125;
                  put_Data_1_1105 <= put_Data_0_1128;
                  put_size_1095 <= put_size_1095 + 1;
                  put_MergeSuccess_1120 <= 1;
                end
                2: begin
                  put_Key_1_1102 <= put_Key_0_1125;
                  put_Data_1_1105 <= put_Data_0_1128;
                  put_Key_2_1106 <= put_Key_1_1129;
                  put_Data_2_1109 <= put_Data_1_1132;
                  put_size_1095 <= put_size_1095 + 2;
                  put_MergeSuccess_1120 <= 1;
                end
                3: begin
                  put_Key_1_1102 <= put_Key_0_1125;
                  put_Data_1_1105 <= put_Data_0_1128;
                  put_Key_2_1106 <= put_Key_1_1129;
                  put_Data_2_1109 <= put_Data_1_1132;
                  put_Key_3_1110 <= put_Key_2_1133;
                  put_Data_3_1113 <= put_Data_2_1136;
                  put_size_1095 <= put_size_1095 + 3;
                  put_MergeSuccess_1120 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1122)
                0: begin
                  put_size_1095 <= put_size_1095 + 0;
                  put_MergeSuccess_1120 <= 1;
                end
                1: begin
                  put_Key_2_1106 <= put_Key_0_1125;
                  put_Data_2_1109 <= put_Data_0_1128;
                  put_size_1095 <= put_size_1095 + 1;
                  put_MergeSuccess_1120 <= 1;
                end
                2: begin
                  put_Key_2_1106 <= put_Key_0_1125;
                  put_Data_2_1109 <= put_Data_0_1128;
                  put_Key_3_1110 <= put_Key_1_1129;
                  put_Data_3_1113 <= put_Data_1_1132;
                  put_size_1095 <= put_size_1095 + 2;
                  put_MergeSuccess_1120 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1122)
                0: begin
                  put_size_1095 <= put_size_1095 + 0;
                  put_MergeSuccess_1120 <= 1;
                end
                1: begin
                  put_Key_3_1110 <= put_Key_0_1125;
                  put_Data_3_1113 <= put_Data_0_1128;
                  put_size_1095 <= put_size_1095 + 1;
                  put_MergeSuccess_1120 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1122)
                0: begin
                  put_size_1095 <= put_size_1095 + 0;
                  put_MergeSuccess_1120 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        701: begin
          if (put_MergeSuccess_1120 == 0) begin
            put_pc <= 724;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        702: begin
          put_size_743 <= put_size_743-1;
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          if (0>= put_StuckIndex_767) begin
            put_Key_0_746 <= put_Key_1_750;
            put_Data_0_749 <= put_Data_1_753;
          end
          if (1>= put_StuckIndex_767) begin
            put_Key_1_750 <= put_Key_2_754;
            put_Data_1_753 <= put_Data_2_757;
          end
          if (2>= put_StuckIndex_767) begin
            put_Key_2_754 <= put_Key_3_758;
            put_Data_2_757 <= put_Data_3_761;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        703: begin
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        704: begin
          if (put_StuckIndex_767 == put_size_743) begin
            put_size_743 <= put_size_743+1;
          end
          case (put_StuckIndex_767)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1150;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1150;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1150;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1150;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        705: begin
          put_success_1153 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        706: begin
          put_stuckSize_6_index_37 <= put_index_1094;
          put_stuckSize_6_value_38 <= put_size_1095;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1094;
          put_stuckKeys_2_value_26 <= put_Key_0_1098;
          put_stuckKeys_2_value_27 <= put_Key_1_1102;
          put_stuckKeys_2_value_28 <= put_Key_2_1106;
          put_stuckKeys_2_value_29 <= put_Key_3_1110;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1094;
          put_stuckData_4_value_32 <= put_Data_0_1101;
          put_stuckData_4_value_33 <= put_Data_1_1105;
          put_stuckData_4_value_34 <= put_Data_2_1109;
          put_stuckData_4_value_35 <= put_Data_3_1113;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        707: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        708: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        709: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        710: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        711: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        712: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        713: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        714: begin
          put_root_1156 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        715: begin
          put_freeNext_9_index_194 <= put_root_1156;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        716: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        717: begin
          put_next_1155 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1156;
          put_freeNext_10_value_196 <= put_indexRight_1151;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1157 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        718: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1151;
          put_stuckIsFree_11_value_198 <= put_isFree_1157;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        719: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        720: begin
          put_freeNext_10_index_195 <= put_indexRight_1151;
          put_freeNext_10_value_196 <= put_next_1155;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        721: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        722: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        723: begin
          put_pc <= 724;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        724: begin
          put_pc <= 725;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        725: begin
          put_pc <= 726;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2470:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        726: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 773;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        727: begin
          put_success_1219 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        728: begin
          case (put_StuckIndex_767)
            0: begin
              put_indexLeft_1216 <= put_Data_0_749;
              put_indexRight_1217 <= put_Data_1_753;
            end
            1: begin
              put_indexLeft_1216 <= put_Data_1_753;
              put_indexRight_1217 <= put_Data_2_757;
            end
            2: begin
              put_indexLeft_1216 <= put_Data_2_757;
              put_indexRight_1217 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        729: begin
          put_index_1158 <= put_indexLeft_1216;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        730: begin
          put_stuckSize_5_index_36 <= put_index_1158;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1158;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1158;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1158;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        731: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        732: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        733: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        734: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        735: begin
          put_size_1159 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1160 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1162 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1165 <= stuckData_stuckData_3_result_0;
          put_Key_1_1166 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1169 <= stuckData_stuckData_3_result_1;
          put_Key_2_1170 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1173 <= stuckData_stuckData_3_result_2;
          put_Key_3_1174 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1177 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        736: begin
          put_index_1185 <= put_indexRight_1217;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        737: begin
          put_stuckSize_5_index_36 <= put_index_1185;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1185;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1185;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1185;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        738: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        739: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        740: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        741: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        742: begin
          put_size_1186 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1187 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1189 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1192 <= stuckData_stuckData_3_result_0;
          put_Key_1_1193 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1196 <= stuckData_stuckData_3_result_1;
          put_Key_2_1197 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1200 <= stuckData_stuckData_3_result_2;
          put_Key_3_1201 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1204 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        743: begin
          if (put_isLeaf_1160 == 0) begin
            put_pc <= 745;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        744: begin
          put_pc <= 773;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        745: begin
          if (put_isLeaf_1187 == 0) begin
            put_pc <= 747;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        746: begin
          put_pc <= 773;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        747: begin
          case (put_StuckIndex_767)
            0: begin
              put_midKey_1218 <= put_Key_0_746;
            end
            1: begin
              put_midKey_1218 <= put_Key_1_750;
            end
            2: begin
              put_midKey_1218 <= put_Key_2_754;
            end
            3: begin
              put_midKey_1218 <= put_Key_3_758;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        748: begin
          put_MergeSuccess_1184 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        749: begin
          case (put_size_1159)
            0: begin
              case (put_size_1186)
                0: begin
                  put_Key_0_1162 <= put_midKey_1218;
                  put_Data_1_1169 <= put_Data_0_1192;
                  put_size_1159 <= put_size_1159 + 1;
                  put_MergeSuccess_1184 <= 1;
                end
                1: begin
                  put_Key_0_1162 <= put_midKey_1218;
                  put_Key_1_1166 <= put_Key_0_1189;
                  put_Data_1_1169 <= put_Data_0_1192;
                  put_Data_2_1173 <= put_Data_1_1196;
                  put_size_1159 <= put_size_1159 + 2;
                  put_MergeSuccess_1184 <= 1;
                end
                2: begin
                  put_Key_0_1162 <= put_midKey_1218;
                  put_Key_1_1166 <= put_Key_0_1189;
                  put_Data_1_1169 <= put_Data_0_1192;
                  put_Key_2_1170 <= put_Key_1_1193;
                  put_Data_2_1173 <= put_Data_1_1196;
                  put_Data_3_1177 <= put_Data_2_1200;
                  put_size_1159 <= put_size_1159 + 3;
                  put_MergeSuccess_1184 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (put_size_1186)
                0: begin
                  put_Key_1_1166 <= put_midKey_1218;
                  put_Data_2_1173 <= put_Data_0_1192;
                  put_size_1159 <= put_size_1159 + 1;
                  put_MergeSuccess_1184 <= 1;
                end
                1: begin
                  put_Key_1_1166 <= put_midKey_1218;
                  put_Key_2_1170 <= put_Key_0_1189;
                  put_Data_2_1173 <= put_Data_0_1192;
                  put_Data_3_1177 <= put_Data_1_1196;
                  put_size_1159 <= put_size_1159 + 2;
                  put_MergeSuccess_1184 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1186)
                0: begin
                  put_Key_2_1170 <= put_midKey_1218;
                  put_Data_3_1177 <= put_Data_0_1192;
                  put_size_1159 <= put_size_1159 + 1;
                  put_MergeSuccess_1184 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1186)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1186)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        750: begin
          if (put_MergeSuccess_1184 == 0) begin
            put_pc <= 773;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        751: begin
          put_size_743 <= put_size_743-1;
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          if (0>= put_StuckIndex_767) begin
            put_Key_0_746 <= put_Key_1_750;
            put_Data_0_749 <= put_Data_1_753;
          end
          if (1>= put_StuckIndex_767) begin
            put_Key_1_750 <= put_Key_2_754;
            put_Data_1_753 <= put_Data_2_757;
          end
          if (2>= put_StuckIndex_767) begin
            put_Key_2_754 <= put_Key_3_758;
            put_Data_2_757 <= put_Data_3_761;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        752: begin
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        753: begin
          if (put_StuckIndex_767 == put_size_743) begin
            put_size_743 <= put_size_743+1;
          end
          case (put_StuckIndex_767)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1216;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1216;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1216;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1216;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        754: begin
          put_success_1219 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        755: begin
          put_stuckSize_6_index_37 <= put_index_1158;
          put_stuckSize_6_value_38 <= put_size_1159;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1158;
          put_stuckKeys_2_value_26 <= put_Key_0_1162;
          put_stuckKeys_2_value_27 <= put_Key_1_1166;
          put_stuckKeys_2_value_28 <= put_Key_2_1170;
          put_stuckKeys_2_value_29 <= put_Key_3_1174;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1158;
          put_stuckData_4_value_32 <= put_Data_0_1165;
          put_stuckData_4_value_33 <= put_Data_1_1169;
          put_stuckData_4_value_34 <= put_Data_2_1173;
          put_stuckData_4_value_35 <= put_Data_3_1177;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        756: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        757: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        758: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        759: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        760: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        761: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        762: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        763: begin
          put_root_1222 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        764: begin
          put_freeNext_9_index_194 <= put_root_1222;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        765: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        766: begin
          put_next_1221 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1222;
          put_freeNext_10_value_196 <= put_indexRight_1217;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1223 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        767: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1217;
          put_stuckIsFree_11_value_198 <= put_isFree_1223;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        768: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        769: begin
          put_freeNext_10_index_195 <= put_indexRight_1217;
          put_freeNext_10_value_196 <= put_next_1221;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        770: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        771: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        772: begin
          put_pc <= 773;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2471:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        773: begin
          put_index1_771 <= put_StuckIndex_767;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2472:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        774: begin
          put_index1_771 <= put_index1_771-1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0813:<init>|  Chip.java:0812:Dec|  Btree.java:2473:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        775: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 819;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        776: begin
          case (put_index1_771)
            0: begin
              put_indexLeft_1280 <= put_Data_0_749;
              put_indexRight_1281 <= put_Data_1_753;
            end
            1: begin
              put_indexLeft_1280 <= put_Data_1_753;
              put_indexRight_1281 <= put_Data_2_757;
            end
            2: begin
              put_indexLeft_1280 <= put_Data_2_757;
              put_indexRight_1281 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        777: begin
          put_index_1224 <= put_indexLeft_1280;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        778: begin
          put_stuckSize_5_index_36 <= put_index_1224;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1224;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1224;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1224;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        779: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        780: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        781: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        782: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        783: begin
          put_size_1225 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1226 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1228 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1231 <= stuckData_stuckData_3_result_0;
          put_Key_1_1232 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1235 <= stuckData_stuckData_3_result_1;
          put_Key_2_1236 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1239 <= stuckData_stuckData_3_result_2;
          put_Key_3_1240 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1243 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        784: begin
          put_index_1251 <= put_indexRight_1281;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        785: begin
          put_stuckSize_5_index_36 <= put_index_1251;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1251;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1251;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1251;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        786: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        787: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        788: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        789: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        790: begin
          put_size_1252 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1253 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1255 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1258 <= stuckData_stuckData_3_result_0;
          put_Key_1_1259 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1262 <= stuckData_stuckData_3_result_1;
          put_Key_2_1263 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1266 <= stuckData_stuckData_3_result_2;
          put_Key_3_1267 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1270 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        791: begin
          if (put_isLeaf_1226 == 0) begin
            put_pc <= 819;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        792: begin
          if (put_isLeaf_1253 == 0) begin
            put_pc <= 818;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        793: begin
          put_MergeSuccess_1250 <= 0;
          case (put_size_1225)
            0: begin
              case (put_size_1252)
                0: begin
                  put_size_1225 <= put_size_1225 + 0;
                  put_MergeSuccess_1250 <= 1;
                end
                1: begin
                  put_Key_0_1228 <= put_Key_0_1255;
                  put_Data_0_1231 <= put_Data_0_1258;
                  put_size_1225 <= put_size_1225 + 1;
                  put_MergeSuccess_1250 <= 1;
                end
                2: begin
                  put_Key_0_1228 <= put_Key_0_1255;
                  put_Data_0_1231 <= put_Data_0_1258;
                  put_Key_1_1232 <= put_Key_1_1259;
                  put_Data_1_1235 <= put_Data_1_1262;
                  put_size_1225 <= put_size_1225 + 2;
                  put_MergeSuccess_1250 <= 1;
                end
                3: begin
                  put_Key_0_1228 <= put_Key_0_1255;
                  put_Data_0_1231 <= put_Data_0_1258;
                  put_Key_1_1232 <= put_Key_1_1259;
                  put_Data_1_1235 <= put_Data_1_1262;
                  put_Key_2_1236 <= put_Key_2_1263;
                  put_Data_2_1239 <= put_Data_2_1266;
                  put_size_1225 <= put_size_1225 + 3;
                  put_MergeSuccess_1250 <= 1;
                end
                4: begin
                  put_Key_0_1228 <= put_Key_0_1255;
                  put_Data_0_1231 <= put_Data_0_1258;
                  put_Key_1_1232 <= put_Key_1_1259;
                  put_Data_1_1235 <= put_Data_1_1262;
                  put_Key_2_1236 <= put_Key_2_1263;
                  put_Data_2_1239 <= put_Data_2_1266;
                  put_Key_3_1240 <= put_Key_3_1267;
                  put_Data_3_1243 <= put_Data_3_1270;
                  put_size_1225 <= put_size_1225 + 4;
                  put_MergeSuccess_1250 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_1252)
                0: begin
                  put_size_1225 <= put_size_1225 + 0;
                  put_MergeSuccess_1250 <= 1;
                end
                1: begin
                  put_Key_1_1232 <= put_Key_0_1255;
                  put_Data_1_1235 <= put_Data_0_1258;
                  put_size_1225 <= put_size_1225 + 1;
                  put_MergeSuccess_1250 <= 1;
                end
                2: begin
                  put_Key_1_1232 <= put_Key_0_1255;
                  put_Data_1_1235 <= put_Data_0_1258;
                  put_Key_2_1236 <= put_Key_1_1259;
                  put_Data_2_1239 <= put_Data_1_1262;
                  put_size_1225 <= put_size_1225 + 2;
                  put_MergeSuccess_1250 <= 1;
                end
                3: begin
                  put_Key_1_1232 <= put_Key_0_1255;
                  put_Data_1_1235 <= put_Data_0_1258;
                  put_Key_2_1236 <= put_Key_1_1259;
                  put_Data_2_1239 <= put_Data_1_1262;
                  put_Key_3_1240 <= put_Key_2_1263;
                  put_Data_3_1243 <= put_Data_2_1266;
                  put_size_1225 <= put_size_1225 + 3;
                  put_MergeSuccess_1250 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1252)
                0: begin
                  put_size_1225 <= put_size_1225 + 0;
                  put_MergeSuccess_1250 <= 1;
                end
                1: begin
                  put_Key_2_1236 <= put_Key_0_1255;
                  put_Data_2_1239 <= put_Data_0_1258;
                  put_size_1225 <= put_size_1225 + 1;
                  put_MergeSuccess_1250 <= 1;
                end
                2: begin
                  put_Key_2_1236 <= put_Key_0_1255;
                  put_Data_2_1239 <= put_Data_0_1258;
                  put_Key_3_1240 <= put_Key_1_1259;
                  put_Data_3_1243 <= put_Data_1_1262;
                  put_size_1225 <= put_size_1225 + 2;
                  put_MergeSuccess_1250 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1252)
                0: begin
                  put_size_1225 <= put_size_1225 + 0;
                  put_MergeSuccess_1250 <= 1;
                end
                1: begin
                  put_Key_3_1240 <= put_Key_0_1255;
                  put_Data_3_1243 <= put_Data_0_1258;
                  put_size_1225 <= put_size_1225 + 1;
                  put_MergeSuccess_1250 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1252)
                0: begin
                  put_size_1225 <= put_size_1225 + 0;
                  put_MergeSuccess_1250 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        794: begin
          if (put_MergeSuccess_1250 == 0) begin
            put_pc <= 817;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        795: begin
          put_size_743 <= put_size_743-1;
          case (put_index1_771)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          if (0>= put_index1_771) begin
            put_Key_0_746 <= put_Key_1_750;
            put_Data_0_749 <= put_Data_1_753;
          end
          if (1>= put_index1_771) begin
            put_Key_1_750 <= put_Key_2_754;
            put_Data_1_753 <= put_Data_2_757;
          end
          if (2>= put_index1_771) begin
            put_Key_2_754 <= put_Key_3_758;
            put_Data_2_757 <= put_Data_3_761;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        796: begin
          case (put_index1_771)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        797: begin
          if (put_index1_771 == put_size_743) begin
            put_size_743 <= put_size_743+1;
          end
          case (put_index1_771)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1280;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1280;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1280;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1280;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        798: begin
          put_success_1283 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        799: begin
          put_stuckSize_6_index_37 <= put_index_1224;
          put_stuckSize_6_value_38 <= put_size_1225;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1224;
          put_stuckKeys_2_value_26 <= put_Key_0_1228;
          put_stuckKeys_2_value_27 <= put_Key_1_1232;
          put_stuckKeys_2_value_28 <= put_Key_2_1236;
          put_stuckKeys_2_value_29 <= put_Key_3_1240;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1224;
          put_stuckData_4_value_32 <= put_Data_0_1231;
          put_stuckData_4_value_33 <= put_Data_1_1235;
          put_stuckData_4_value_34 <= put_Data_2_1239;
          put_stuckData_4_value_35 <= put_Data_3_1243;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        800: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        801: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        802: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        803: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        804: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        805: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        806: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        807: begin
          put_root_1286 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        808: begin
          put_freeNext_9_index_194 <= put_root_1286;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        809: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        810: begin
          put_next_1285 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1286;
          put_freeNext_10_value_196 <= put_indexRight_1281;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1287 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        811: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1281;
          put_stuckIsFree_11_value_198 <= put_isFree_1287;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        812: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        813: begin
          put_freeNext_10_index_195 <= put_indexRight_1281;
          put_freeNext_10_value_196 <= put_next_1285;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        814: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        815: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        816: begin
          put_pc <= 817;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        817: begin
          put_pc <= 818;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        818: begin
          put_pc <= 819;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2474:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        819: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 866;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        820: begin
          put_success_1349 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        821: begin
          case (put_index1_771)
            0: begin
              put_indexLeft_1346 <= put_Data_0_749;
              put_indexRight_1347 <= put_Data_1_753;
            end
            1: begin
              put_indexLeft_1346 <= put_Data_1_753;
              put_indexRight_1347 <= put_Data_2_757;
            end
            2: begin
              put_indexLeft_1346 <= put_Data_2_757;
              put_indexRight_1347 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        822: begin
          put_index_1288 <= put_indexLeft_1346;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        823: begin
          put_stuckSize_5_index_36 <= put_index_1288;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1288;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1288;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1288;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        824: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        825: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        826: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        827: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        828: begin
          put_size_1289 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1290 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1292 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1295 <= stuckData_stuckData_3_result_0;
          put_Key_1_1296 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1299 <= stuckData_stuckData_3_result_1;
          put_Key_2_1300 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1303 <= stuckData_stuckData_3_result_2;
          put_Key_3_1304 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1307 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        829: begin
          put_index_1315 <= put_indexRight_1347;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        830: begin
          put_stuckSize_5_index_36 <= put_index_1315;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1315;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1315;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1315;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        831: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        832: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        833: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        834: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        835: begin
          put_size_1316 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1317 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1319 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1322 <= stuckData_stuckData_3_result_0;
          put_Key_1_1323 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1326 <= stuckData_stuckData_3_result_1;
          put_Key_2_1327 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1330 <= stuckData_stuckData_3_result_2;
          put_Key_3_1331 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1334 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        836: begin
          if (put_isLeaf_1290 == 0) begin
            put_pc <= 838;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        837: begin
          put_pc <= 866;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        838: begin
          if (put_isLeaf_1317 == 0) begin
            put_pc <= 840;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        839: begin
          put_pc <= 866;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        840: begin
          case (put_index1_771)
            0: begin
              put_midKey_1348 <= put_Key_0_746;
            end
            1: begin
              put_midKey_1348 <= put_Key_1_750;
            end
            2: begin
              put_midKey_1348 <= put_Key_2_754;
            end
            3: begin
              put_midKey_1348 <= put_Key_3_758;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        841: begin
          put_MergeSuccess_1314 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        842: begin
          case (put_size_1289)
            0: begin
              case (put_size_1316)
                0: begin
                  put_Key_0_1292 <= put_midKey_1348;
                  put_Data_1_1299 <= put_Data_0_1322;
                  put_size_1289 <= put_size_1289 + 1;
                  put_MergeSuccess_1314 <= 1;
                end
                1: begin
                  put_Key_0_1292 <= put_midKey_1348;
                  put_Key_1_1296 <= put_Key_0_1319;
                  put_Data_1_1299 <= put_Data_0_1322;
                  put_Data_2_1303 <= put_Data_1_1326;
                  put_size_1289 <= put_size_1289 + 2;
                  put_MergeSuccess_1314 <= 1;
                end
                2: begin
                  put_Key_0_1292 <= put_midKey_1348;
                  put_Key_1_1296 <= put_Key_0_1319;
                  put_Data_1_1299 <= put_Data_0_1322;
                  put_Key_2_1300 <= put_Key_1_1323;
                  put_Data_2_1303 <= put_Data_1_1326;
                  put_Data_3_1307 <= put_Data_2_1330;
                  put_size_1289 <= put_size_1289 + 3;
                  put_MergeSuccess_1314 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (put_size_1316)
                0: begin
                  put_Key_1_1296 <= put_midKey_1348;
                  put_Data_2_1303 <= put_Data_0_1322;
                  put_size_1289 <= put_size_1289 + 1;
                  put_MergeSuccess_1314 <= 1;
                end
                1: begin
                  put_Key_1_1296 <= put_midKey_1348;
                  put_Key_2_1300 <= put_Key_0_1319;
                  put_Data_2_1303 <= put_Data_0_1322;
                  put_Data_3_1307 <= put_Data_1_1326;
                  put_size_1289 <= put_size_1289 + 2;
                  put_MergeSuccess_1314 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1316)
                0: begin
                  put_Key_2_1300 <= put_midKey_1348;
                  put_Data_3_1307 <= put_Data_0_1322;
                  put_size_1289 <= put_size_1289 + 1;
                  put_MergeSuccess_1314 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1316)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1316)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        843: begin
          if (put_MergeSuccess_1314 == 0) begin
            put_pc <= 866;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        844: begin
          put_size_743 <= put_size_743-1;
          case (put_index1_771)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          if (0>= put_index1_771) begin
            put_Key_0_746 <= put_Key_1_750;
            put_Data_0_749 <= put_Data_1_753;
          end
          if (1>= put_index1_771) begin
            put_Key_1_750 <= put_Key_2_754;
            put_Data_1_753 <= put_Data_2_757;
          end
          if (2>= put_index1_771) begin
            put_Key_2_754 <= put_Key_3_758;
            put_Data_2_757 <= put_Data_3_761;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        845: begin
          case (put_index1_771)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        846: begin
          if (put_index1_771 == put_size_743) begin
            put_size_743 <= put_size_743+1;
          end
          case (put_index1_771)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1346;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1346;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1346;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1346;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        847: begin
          put_success_1349 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        848: begin
          put_stuckSize_6_index_37 <= put_index_1288;
          put_stuckSize_6_value_38 <= put_size_1289;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1288;
          put_stuckKeys_2_value_26 <= put_Key_0_1292;
          put_stuckKeys_2_value_27 <= put_Key_1_1296;
          put_stuckKeys_2_value_28 <= put_Key_2_1300;
          put_stuckKeys_2_value_29 <= put_Key_3_1304;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1288;
          put_stuckData_4_value_32 <= put_Data_0_1295;
          put_stuckData_4_value_33 <= put_Data_1_1299;
          put_stuckData_4_value_34 <= put_Data_2_1303;
          put_stuckData_4_value_35 <= put_Data_3_1307;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        849: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        850: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        851: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        852: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        853: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        854: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        855: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        856: begin
          put_root_1352 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        857: begin
          put_freeNext_9_index_194 <= put_root_1352;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        858: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        859: begin
          put_next_1351 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1352;
          put_freeNext_10_value_196 <= put_indexRight_1347;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1353 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        860: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1347;
          put_stuckIsFree_11_value_198 <= put_isFree_1353;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        861: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        862: begin
          put_freeNext_10_index_195 <= put_indexRight_1347;
          put_freeNext_10_value_196 <= put_next_1351;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        863: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        864: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        865: begin
          put_pc <= 866;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2475:Then|  Chip.java:0610:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        866: begin
          put_pc <= 958;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        867: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 911;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:1876:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        868: begin
          case (put_StuckIndex_767)
            0: begin
              put_indexLeft_1410 <= put_Data_0_749;
              put_indexRight_1411 <= put_Data_1_753;
            end
            1: begin
              put_indexLeft_1410 <= put_Data_1_753;
              put_indexRight_1411 <= put_Data_2_757;
            end
            2: begin
              put_indexLeft_1410 <= put_Data_2_757;
              put_indexRight_1411 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1879:<init>|  Btree.java:1878:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        869: begin
          put_index_1354 <= put_indexLeft_1410;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        870: begin
          put_stuckSize_5_index_36 <= put_index_1354;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1354;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1354;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1354;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        871: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        872: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        873: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        874: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        875: begin
          put_size_1355 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1356 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1358 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1361 <= stuckData_stuckData_3_result_0;
          put_Key_1_1362 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1365 <= stuckData_stuckData_3_result_1;
          put_Key_2_1366 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1369 <= stuckData_stuckData_3_result_2;
          put_Key_3_1370 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1373 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1893:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        876: begin
          put_index_1381 <= put_indexRight_1411;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        877: begin
          put_stuckSize_5_index_36 <= put_index_1381;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1381;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1381;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1381;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        878: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        879: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        880: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        881: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        882: begin
          put_size_1382 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1383 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1385 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1388 <= stuckData_stuckData_3_result_0;
          put_Key_1_1389 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1392 <= stuckData_stuckData_3_result_1;
          put_Key_2_1393 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1396 <= stuckData_stuckData_3_result_2;
          put_Key_3_1397 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1400 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:1894:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        883: begin
          if (put_isLeaf_1356 == 0) begin
            put_pc <= 911;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        884: begin
          if (put_isLeaf_1383 == 0) begin
            put_pc <= 910;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        885: begin
          put_MergeSuccess_1380 <= 0;
          case (put_size_1355)
            0: begin
              case (put_size_1382)
                0: begin
                  put_size_1355 <= put_size_1355 + 0;
                  put_MergeSuccess_1380 <= 1;
                end
                1: begin
                  put_Key_0_1358 <= put_Key_0_1385;
                  put_Data_0_1361 <= put_Data_0_1388;
                  put_size_1355 <= put_size_1355 + 1;
                  put_MergeSuccess_1380 <= 1;
                end
                2: begin
                  put_Key_0_1358 <= put_Key_0_1385;
                  put_Data_0_1361 <= put_Data_0_1388;
                  put_Key_1_1362 <= put_Key_1_1389;
                  put_Data_1_1365 <= put_Data_1_1392;
                  put_size_1355 <= put_size_1355 + 2;
                  put_MergeSuccess_1380 <= 1;
                end
                3: begin
                  put_Key_0_1358 <= put_Key_0_1385;
                  put_Data_0_1361 <= put_Data_0_1388;
                  put_Key_1_1362 <= put_Key_1_1389;
                  put_Data_1_1365 <= put_Data_1_1392;
                  put_Key_2_1366 <= put_Key_2_1393;
                  put_Data_2_1369 <= put_Data_2_1396;
                  put_size_1355 <= put_size_1355 + 3;
                  put_MergeSuccess_1380 <= 1;
                end
                4: begin
                  put_Key_0_1358 <= put_Key_0_1385;
                  put_Data_0_1361 <= put_Data_0_1388;
                  put_Key_1_1362 <= put_Key_1_1389;
                  put_Data_1_1365 <= put_Data_1_1392;
                  put_Key_2_1366 <= put_Key_2_1393;
                  put_Data_2_1369 <= put_Data_2_1396;
                  put_Key_3_1370 <= put_Key_3_1397;
                  put_Data_3_1373 <= put_Data_3_1400;
                  put_size_1355 <= put_size_1355 + 4;
                  put_MergeSuccess_1380 <= 1;
                end
              endcase
            end
            1: begin
              case (put_size_1382)
                0: begin
                  put_size_1355 <= put_size_1355 + 0;
                  put_MergeSuccess_1380 <= 1;
                end
                1: begin
                  put_Key_1_1362 <= put_Key_0_1385;
                  put_Data_1_1365 <= put_Data_0_1388;
                  put_size_1355 <= put_size_1355 + 1;
                  put_MergeSuccess_1380 <= 1;
                end
                2: begin
                  put_Key_1_1362 <= put_Key_0_1385;
                  put_Data_1_1365 <= put_Data_0_1388;
                  put_Key_2_1366 <= put_Key_1_1389;
                  put_Data_2_1369 <= put_Data_1_1392;
                  put_size_1355 <= put_size_1355 + 2;
                  put_MergeSuccess_1380 <= 1;
                end
                3: begin
                  put_Key_1_1362 <= put_Key_0_1385;
                  put_Data_1_1365 <= put_Data_0_1388;
                  put_Key_2_1366 <= put_Key_1_1389;
                  put_Data_2_1369 <= put_Data_1_1392;
                  put_Key_3_1370 <= put_Key_2_1393;
                  put_Data_3_1373 <= put_Data_2_1396;
                  put_size_1355 <= put_size_1355 + 3;
                  put_MergeSuccess_1380 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1382)
                0: begin
                  put_size_1355 <= put_size_1355 + 0;
                  put_MergeSuccess_1380 <= 1;
                end
                1: begin
                  put_Key_2_1366 <= put_Key_0_1385;
                  put_Data_2_1369 <= put_Data_0_1388;
                  put_size_1355 <= put_size_1355 + 1;
                  put_MergeSuccess_1380 <= 1;
                end
                2: begin
                  put_Key_2_1366 <= put_Key_0_1385;
                  put_Data_2_1369 <= put_Data_0_1388;
                  put_Key_3_1370 <= put_Key_1_1389;
                  put_Data_3_1373 <= put_Data_1_1392;
                  put_size_1355 <= put_size_1355 + 2;
                  put_MergeSuccess_1380 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1382)
                0: begin
                  put_size_1355 <= put_size_1355 + 0;
                  put_MergeSuccess_1380 <= 1;
                end
                1: begin
                  put_Key_3_1370 <= put_Key_0_1385;
                  put_Data_3_1373 <= put_Data_0_1388;
                  put_size_1355 <= put_size_1355 + 1;
                  put_MergeSuccess_1380 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1382)
                0: begin
                  put_size_1355 <= put_size_1355 + 0;
                  put_MergeSuccess_1380 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1212:<init>|  Btree.java:1211:merge|  Btree.java:1900:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        886: begin
          if (put_MergeSuccess_1380 == 0) begin
            put_pc <= 909;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        887: begin
          put_size_743 <= put_size_743-1;
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          if (0>= put_StuckIndex_767) begin
            put_Key_0_746 <= put_Key_1_750;
            put_Data_0_749 <= put_Data_1_753;
          end
          if (1>= put_StuckIndex_767) begin
            put_Key_1_750 <= put_Key_2_754;
            put_Data_1_753 <= put_Data_2_757;
          end
          if (2>= put_StuckIndex_767) begin
            put_Key_2_754 <= put_Key_3_758;
            put_Data_2_757 <= put_Data_3_761;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:1904:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        888: begin
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:1905:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        889: begin
          if (put_StuckIndex_767 == put_size_743) begin
            put_size_743 <= put_size_743+1;
          end
          case (put_StuckIndex_767)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1410;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1410;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1410;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1410;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:1906:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        890: begin
          put_success_1413 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:1907:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        891: begin
          put_stuckSize_6_index_37 <= put_index_1354;
          put_stuckSize_6_value_38 <= put_size_1355;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1354;
          put_stuckKeys_2_value_26 <= put_Key_0_1358;
          put_stuckKeys_2_value_27 <= put_Key_1_1362;
          put_stuckKeys_2_value_28 <= put_Key_2_1366;
          put_stuckKeys_2_value_29 <= put_Key_3_1370;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1354;
          put_stuckData_4_value_32 <= put_Data_0_1361;
          put_stuckData_4_value_33 <= put_Data_1_1365;
          put_stuckData_4_value_34 <= put_Data_2_1369;
          put_stuckData_4_value_35 <= put_Data_3_1373;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        892: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        893: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        894: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1908:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        895: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        896: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        897: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        898: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:1909:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        899: begin
          put_root_1416 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        900: begin
          put_freeNext_9_index_194 <= put_root_1416;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        901: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        902: begin
          put_next_1415 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1416;
          put_freeNext_10_value_196 <= put_indexRight_1411;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1417 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        903: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1411;
          put_stuckIsFree_11_value_198 <= put_isFree_1417;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        904: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        905: begin
          put_freeNext_10_index_195 <= put_indexRight_1411;
          put_freeNext_10_value_196 <= put_next_1415;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        906: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        907: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:1910:Then|  Chip.java:0610:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        908: begin
          put_pc <= 909;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:1903:<init>|  Btree.java:1902:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        909: begin
          put_pc <= 910;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1899:<init>|  Btree.java:1898:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        910: begin
          put_pc <= 911;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:1897:<init>|  Btree.java:1896:code|  Chip.java:0530:<init>|  Btree.java:1875:<init>|  Btree.java:1874:mergeLeavesNotTop|  Btree.java:2478:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        911: begin
          if (put_position_769 == 0 && put_size_743 > 1) begin
            put_pc <= put_pc + 1;
          end
          else begin
            if (put_position_769 == 0 || put_size_743 < 1) begin
              put_pc <= 958;
            end
            else begin
              put_pc <= put_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2100:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        912: begin
          put_success_1479 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2101:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        913: begin
          case (put_StuckIndex_767)
            0: begin
              put_indexLeft_1476 <= put_Data_0_749;
              put_indexRight_1477 <= put_Data_1_753;
            end
            1: begin
              put_indexLeft_1476 <= put_Data_1_753;
              put_indexRight_1477 <= put_Data_2_757;
            end
            2: begin
              put_indexLeft_1476 <= put_Data_2_757;
              put_indexRight_1477 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2104:<init>|  Btree.java:2103:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        914: begin
          put_index_1418 <= put_indexLeft_1476;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        915: begin
          put_stuckSize_5_index_36 <= put_index_1418;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1418;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1418;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1418;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        916: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        917: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        918: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        919: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        920: begin
          put_size_1419 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1420 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1422 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1425 <= stuckData_stuckData_3_result_0;
          put_Key_1_1426 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1429 <= stuckData_stuckData_3_result_1;
          put_Key_2_1430 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1433 <= stuckData_stuckData_3_result_2;
          put_Key_3_1434 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1437 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2118:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        921: begin
          put_index_1445 <= put_indexRight_1477;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        922: begin
          put_stuckSize_5_index_36 <= put_index_1445;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_1445;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_1445;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_1445;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        923: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        924: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        925: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        926: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        927: begin
          put_size_1446 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_1447 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_1449 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_1452 <= stuckData_stuckData_3_result_0;
          put_Key_1_1453 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_1456 <= stuckData_stuckData_3_result_1;
          put_Key_2_1457 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_1460 <= stuckData_stuckData_3_result_2;
          put_Key_3_1461 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_1464 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2119:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        928: begin
          if (put_isLeaf_1420 == 0) begin
            put_pc <= 930;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        929: begin
          put_pc <= 958;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        930: begin
          if (put_isLeaf_1447 == 0) begin
            put_pc <= 932;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        931: begin
          put_pc <= 958;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        932: begin
          case (put_StuckIndex_767)
            0: begin
              put_midKey_1478 <= put_Key_0_746;
            end
            1: begin
              put_midKey_1478 <= put_Key_1_750;
            end
            2: begin
              put_midKey_1478 <= put_Key_2_754;
            end
            3: begin
              put_midKey_1478 <= put_Key_3_758;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2126:<init>|  Btree.java:2125:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        933: begin
          put_MergeSuccess_1444 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        934: begin
          case (put_size_1419)
            0: begin
              case (put_size_1446)
                0: begin
                  put_Key_0_1422 <= put_midKey_1478;
                  put_Data_1_1429 <= put_Data_0_1452;
                  put_size_1419 <= put_size_1419 + 1;
                  put_MergeSuccess_1444 <= 1;
                end
                1: begin
                  put_Key_0_1422 <= put_midKey_1478;
                  put_Key_1_1426 <= put_Key_0_1449;
                  put_Data_1_1429 <= put_Data_0_1452;
                  put_Data_2_1433 <= put_Data_1_1456;
                  put_size_1419 <= put_size_1419 + 2;
                  put_MergeSuccess_1444 <= 1;
                end
                2: begin
                  put_Key_0_1422 <= put_midKey_1478;
                  put_Key_1_1426 <= put_Key_0_1449;
                  put_Data_1_1429 <= put_Data_0_1452;
                  put_Key_2_1430 <= put_Key_1_1453;
                  put_Data_2_1433 <= put_Data_1_1456;
                  put_Data_3_1437 <= put_Data_2_1460;
                  put_size_1419 <= put_size_1419 + 3;
                  put_MergeSuccess_1444 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (put_size_1446)
                0: begin
                  put_Key_1_1426 <= put_midKey_1478;
                  put_Data_2_1433 <= put_Data_0_1452;
                  put_size_1419 <= put_size_1419 + 1;
                  put_MergeSuccess_1444 <= 1;
                end
                1: begin
                  put_Key_1_1426 <= put_midKey_1478;
                  put_Key_2_1430 <= put_Key_0_1449;
                  put_Data_2_1433 <= put_Data_0_1452;
                  put_Data_3_1437 <= put_Data_1_1456;
                  put_size_1419 <= put_size_1419 + 2;
                  put_MergeSuccess_1444 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (put_size_1446)
                0: begin
                  put_Key_2_1430 <= put_midKey_1478;
                  put_Data_3_1437 <= put_Data_0_1452;
                  put_size_1419 <= put_size_1419 + 1;
                  put_MergeSuccess_1444 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (put_size_1446)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (put_size_1446)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2138:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        935: begin
          if (put_MergeSuccess_1444 == 0) begin
            put_pc <= 958;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        936: begin
          put_size_743 <= put_size_743-1;
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          if (0>= put_StuckIndex_767) begin
            put_Key_0_746 <= put_Key_1_750;
            put_Data_0_749 <= put_Data_1_753;
          end
          if (1>= put_StuckIndex_767) begin
            put_Key_1_750 <= put_Key_2_754;
            put_Data_1_753 <= put_Data_2_757;
          end
          if (2>= put_StuckIndex_767) begin
            put_Key_2_754 <= put_Key_3_758;
            put_Data_2_757 <= put_Data_3_761;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0742:<init>|  Btree.java:0741:RemoveElementAt|  Btree.java:2142:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        937: begin
          case (put_StuckIndex_767)
            0: begin
              put_Key_763 <= put_Key_0_746;
              put_Data_765 <= put_Data_0_749;
            end
            1: begin
              put_Key_763 <= put_Key_1_750;
              put_Data_765 <= put_Data_1_753;
            end
            2: begin
              put_Key_763 <= put_Key_2_754;
              put_Data_765 <= put_Data_2_757;
            end
            3: begin
              put_Key_763 <= put_Key_3_758;
              put_Data_765 <= put_Data_3_761;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0583:<init>|  Btree.java:0582:ElementAt|  Btree.java:2143:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        938: begin
          if (put_StuckIndex_767 == put_size_743) begin
            put_size_743 <= put_size_743+1;
          end
          case (put_StuckIndex_767)
            0: begin
              put_Key_0_746 <= put_Key_763;
              put_Data_0_749 <= put_indexLeft_1476;
            end
            1: begin
              put_Key_1_750 <= put_Key_763;
              put_Data_1_753 <= put_indexLeft_1476;
            end
            2: begin
              put_Key_2_754 <= put_Key_763;
              put_Data_2_757 <= put_indexLeft_1476;
            end
            3: begin
              put_Key_3_758 <= put_Key_763;
              put_Data_3_761 <= put_indexLeft_1476;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0625:<init>|  Btree.java:0624:SetElementAt|  Btree.java:2144:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        939: begin
          put_success_1479 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2145:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        940: begin
          put_stuckSize_6_index_37 <= put_index_1418;
          put_stuckSize_6_value_38 <= put_size_1419;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_1418;
          put_stuckKeys_2_value_26 <= put_Key_0_1422;
          put_stuckKeys_2_value_27 <= put_Key_1_1426;
          put_stuckKeys_2_value_28 <= put_Key_2_1430;
          put_stuckKeys_2_value_29 <= put_Key_3_1434;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_1418;
          put_stuckData_4_value_32 <= put_Data_0_1425;
          put_stuckData_4_value_33 <= put_Data_1_1429;
          put_stuckData_4_value_34 <= put_Data_2_1433;
          put_stuckData_4_value_35 <= put_Data_3_1437;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        941: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        942: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        943: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2146:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        944: begin
          put_stuckSize_6_index_37 <= put_index_742;
          put_stuckSize_6_value_38 <= put_size_743;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_742;
          put_stuckKeys_2_value_26 <= put_Key_0_746;
          put_stuckKeys_2_value_27 <= put_Key_1_750;
          put_stuckKeys_2_value_28 <= put_Key_2_754;
          put_stuckKeys_2_value_29 <= put_Key_3_758;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_742;
          put_stuckData_4_value_32 <= put_Data_0_749;
          put_stuckData_4_value_33 <= put_Data_1_753;
          put_stuckData_4_value_34 <= put_Data_2_757;
          put_stuckData_4_value_35 <= put_Data_3_761;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        945: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        946: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        947: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2147:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        948: begin
          put_root_1482 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        949: begin
          put_freeNext_9_index_194 <= put_root_1482;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        950: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        951: begin
          put_next_1481 <= freeNext_freeNext_9_result_0;
          put_freeNext_10_index_195 <= put_root_1482;
          put_freeNext_10_value_196 <= put_indexRight_1477;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_isFree_1483 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        952: begin
          put_stuckIsFree_11_index_197 <= put_indexRight_1477;
          put_stuckIsFree_11_value_198 <= put_isFree_1483;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        953: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        954: begin
          put_freeNext_10_index_195 <= put_indexRight_1477;
          put_freeNext_10_value_196 <= put_next_1481;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        955: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        956: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2148:Then|  Chip.java:0610:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        957: begin
          put_pc <= 958;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2141:<init>|  Btree.java:2140:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2124:<init>|  Btree.java:2123:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2122:<init>|  Btree.java:2121:code|  Chip.java:0530:<init>|  Btree.java:2099:<init>|  Btree.java:2098:mergeBranchesNotTop|  Btree.java:2479:Else|  Chip.java:0620:<init>|  Btree.java:2469:<init>|  Btree.java:2468:Then|  Chip.java:0610:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        958: begin
          put_pc <= 959;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2467:<init>|  Btree.java:2466:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        959: begin
          put_index_742 <= put_position_769;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        960: begin
          put_stuckSize_5_index_36 <= put_index_742;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_742;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_742;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_742;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        961: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        962: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        963: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        964: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        965: begin
          put_size_743 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_744 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_746 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_749 <= stuckData_stuckData_3_result_0;
          put_Key_1_750 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_753 <= stuckData_stuckData_3_result_1;
          put_Key_2_754 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_757 <= stuckData_stuckData_3_result_2;
          put_Key_3_758 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_761 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2485:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        966: begin
          put_KeyCompares_0_747 <= put_k_0 <= put_Key_0_746 && 0 < put_size_743;
          put_KeyCollapse_0_748 <= 0;
          put_KeyCompares_1_751 <= put_k_0 >  put_Key_0_746 && put_k_0 <= put_Key_1_750 && 1 < put_size_743;
          put_KeyCollapse_1_752 <= 1;
          put_KeyCompares_2_755 <= put_k_0 >  put_Key_1_750 && put_k_0 <= put_Key_2_754 && 2 < put_size_743;
          put_KeyCollapse_2_756 <= 2;
          put_KeyCompares_3_759 <= put_k_0 >  put_Key_2_754 && put_k_0 <= put_Key_3_758 && 3 < put_size_743;
          put_KeyCollapse_3_760 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0937:<init>|  Btree.java:0936:search_le_parallel|  Btree.java:2487:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        967: begin
          if (put_KeyCompares_1_751) begin
            put_KeyCompares_0_747 <= 1;
            put_KeyCollapse_0_748 <= put_KeyCollapse_1_752;
          end
          if (put_KeyCompares_3_759) begin
            put_KeyCompares_2_755 <= 1;
            put_KeyCollapse_2_756 <= put_KeyCollapse_3_760;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2487:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        968: begin
          if (put_KeyCompares_2_755) begin
            put_KeyCompares_0_747 <= 1;
            put_KeyCollapse_0_748 <= put_KeyCollapse_2_756;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0973:<init>|  Btree.java:0972:search_le_parallel|  Btree.java:2487:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        969: begin
          if (put_KeyCompares_0_747) begin
            put_Found_762 <= 1;
            case (put_KeyCollapse_0_748)
              0: begin
                put_StuckIndex_767 <= 0;
                put_FoundKey_764 <= put_Key_0_746;
                put_Data_765 <= put_Data_0_749;
              end
              1: begin
                put_StuckIndex_767 <= 1;
                put_FoundKey_764 <= put_Key_1_750;
                put_Data_765 <= put_Data_1_753;
              end
              2: begin
                put_StuckIndex_767 <= 2;
                put_FoundKey_764 <= put_Key_2_754;
                put_Data_765 <= put_Data_2_757;
              end
              3: begin
                put_StuckIndex_767 <= 3;
                put_FoundKey_764 <= put_Key_3_758;
                put_Data_765 <= put_Data_3_761;
              end
            endcase
          end
          else begin
            put_Found_762 <= 0;
            case (put_size_743)
              0: begin
                put_StuckIndex_767 <= 0;
                put_Data_765 <= put_Data_0_749;
              end
              1: begin
                put_StuckIndex_767 <= 1;
                put_Data_765 <= put_Data_1_753;
              end
              2: begin
                put_StuckIndex_767 <= 2;
                put_Data_765 <= put_Data_2_757;
              end
              3: begin
                put_StuckIndex_767 <= 3;
                put_Data_765 <= put_Data_3_761;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0995:<init>|  Btree.java:0994:search_le_parallel|  Btree.java:2487:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        970: begin
          put_position_769 <= put_Data_765;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2488:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        971: begin
          put_index_742 <= put_position_769;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        972: begin
          put_stuckSize_5_index_36 <= put_index_742;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_742;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_742;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_742;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        973: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        974: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        975: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        976: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        977: begin
          put_size_743 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_744 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_746 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_749 <= stuckData_stuckData_3_result_0;
          put_Key_1_750 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_753 <= stuckData_stuckData_3_result_1;
          put_Key_2_754 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_757 <= stuckData_stuckData_3_result_2;
          put_Key_3_758 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_761 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2490:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        978: begin
          if (put_isLeaf_744 == 0) begin
            put_pc <= 981;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2493:<init>|  Btree.java:2492:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        979: begin
          put_pc <= 982;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2494:Leaf|  Btree.java:1409:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2493:<init>|  Btree.java:2492:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        980: begin
          put_pc <= 982;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2493:<init>|  Btree.java:2492:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        981: begin
          put_pc <= 587;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2497:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2493:<init>|  Btree.java:2492:code|  Chip.java:0530:<init>|  Btree.java:2456:<init>|  Btree.java:2455:code|  Chip.java:0530:<init>|  Btree.java:2433:<init>|  Btree.java:2432:merge|  Btree.java:2420:put|  Btree.java:6069:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        982: begin
          put_l_3 <= put_k_0< 32 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:6071:<init>|  Btree.java:6070:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        983: begin
          if (put_l_3 >  0) begin
            put_pc <= 0;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0578:<init>|  Chip.java:0577:GONotZero|  Btree.java:6079:code|  Chip.java:0530:<init>|  Btree.java:6067:<init>|  Btree.java:6066:test_put_merge|  Btree.java:7012:newTests|  Btree.java:7018:main|");
            $fclose(f);
          end
        end
        default: put_stop <= 1;
      endcase
    end
  end
  task chipPrint;
    begin
      integer o;
      o = $fopen("verilog/trace_verilog.txt", "a");
      if (!o) o = $fopen("../verilog/trace_verilog.txt", "a");
      if (!o) $display("Cannot create trace folder: verilog/trace_verilog.txt");
      $fwrite(o, "Chip: %-16s step: %1d, maxSteps: %1d, running: %1d\n", "Btree", step, maxSteps, !stop);
      $fwrite(o, "  Processes:\n");

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 0, "stuckIsLeaf", 1, stuckIsLeaf_pc, stuckIsLeaf_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsLeaf_memory[0]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[1]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[2]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[3]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[4]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[5]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[6]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[7]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[8]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[9]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[10]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[11]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[12]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[13]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[14]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[15]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[16]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[17]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[18]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[19]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[20]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[21]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[22]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[23]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[24]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[25]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[26]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[27]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[28]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[29]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[30]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckIsLeaf_7", stuckIsLeaf_7_requestedAt, stuckIsLeaf_7_finishedAt, stuckIsLeaf_stuckIsLeaf_7_returnCode, (stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step), (stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsLeaf_7_index_39", put_stuckIsLeaf_7_index_39);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsLeaf_8", stuckIsLeaf_8_requestedAt, stuckIsLeaf_8_finishedAt, stuckIsLeaf_stuckIsLeaf_8_returnCode, (stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step), (stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsLeaf_8_index_40", put_stuckIsLeaf_8_index_40);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsLeaf_8_value_41", put_stuckIsLeaf_8_value_41);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 1, "stuckIsFree", 1, stuckIsFree_pc, stuckIsFree_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsFree_memory[0]);
      $fwrite(o, ", %2d", stuckIsFree_memory[1]);
      $fwrite(o, ", %2d", stuckIsFree_memory[2]);
      $fwrite(o, ", %2d", stuckIsFree_memory[3]);
      $fwrite(o, ", %2d", stuckIsFree_memory[4]);
      $fwrite(o, ", %2d", stuckIsFree_memory[5]);
      $fwrite(o, ", %2d", stuckIsFree_memory[6]);
      $fwrite(o, ", %2d", stuckIsFree_memory[7]);
      $fwrite(o, ", %2d", stuckIsFree_memory[8]);
      $fwrite(o, ", %2d", stuckIsFree_memory[9]);
      $fwrite(o, ", %2d", stuckIsFree_memory[10]);
      $fwrite(o, ", %2d", stuckIsFree_memory[11]);
      $fwrite(o, ", %2d", stuckIsFree_memory[12]);
      $fwrite(o, ", %2d", stuckIsFree_memory[13]);
      $fwrite(o, ", %2d", stuckIsFree_memory[14]);
      $fwrite(o, ", %2d", stuckIsFree_memory[15]);
      $fwrite(o, ", %2d", stuckIsFree_memory[16]);
      $fwrite(o, ", %2d", stuckIsFree_memory[17]);
      $fwrite(o, ", %2d", stuckIsFree_memory[18]);
      $fwrite(o, ", %2d", stuckIsFree_memory[19]);
      $fwrite(o, ", %2d", stuckIsFree_memory[20]);
      $fwrite(o, ", %2d", stuckIsFree_memory[21]);
      $fwrite(o, ", %2d", stuckIsFree_memory[22]);
      $fwrite(o, ", %2d", stuckIsFree_memory[23]);
      $fwrite(o, ", %2d", stuckIsFree_memory[24]);
      $fwrite(o, ", %2d", stuckIsFree_memory[25]);
      $fwrite(o, ", %2d", stuckIsFree_memory[26]);
      $fwrite(o, ", %2d", stuckIsFree_memory[27]);
      $fwrite(o, ", %2d", stuckIsFree_memory[28]);
      $fwrite(o, ", %2d", stuckIsFree_memory[29]);
      $fwrite(o, ", %2d", stuckIsFree_memory[30]);
      $fwrite(o, ", %2d", stuckIsFree_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsFree_11", stuckIsFree_11_requestedAt, stuckIsFree_11_finishedAt, stuckIsFree_stuckIsFree_11_returnCode, (stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step), (stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsFree_11_index_197", put_stuckIsFree_11_index_197);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsFree_11_value_198", put_stuckIsFree_11_value_198);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 2, "freeNext", 1, freeNext_pc, freeNext_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 6, 1);
      $fwrite(o, "        %2d", freeNext_memory[0]);
      $fwrite(o, ", %2d", freeNext_memory[1]);
      $fwrite(o, ", %2d", freeNext_memory[2]);
      $fwrite(o, ", %2d", freeNext_memory[3]);
      $fwrite(o, ", %2d", freeNext_memory[4]);
      $fwrite(o, ", %2d", freeNext_memory[5]);
      $fwrite(o, ", %2d", freeNext_memory[6]);
      $fwrite(o, ", %2d", freeNext_memory[7]);
      $fwrite(o, ", %2d", freeNext_memory[8]);
      $fwrite(o, ", %2d", freeNext_memory[9]);
      $fwrite(o, ", %2d", freeNext_memory[10]);
      $fwrite(o, ", %2d", freeNext_memory[11]);
      $fwrite(o, ", %2d", freeNext_memory[12]);
      $fwrite(o, ", %2d", freeNext_memory[13]);
      $fwrite(o, ", %2d", freeNext_memory[14]);
      $fwrite(o, ", %2d", freeNext_memory[15]);
      $fwrite(o, ", %2d", freeNext_memory[16]);
      $fwrite(o, ", %2d", freeNext_memory[17]);
      $fwrite(o, ", %2d", freeNext_memory[18]);
      $fwrite(o, ", %2d", freeNext_memory[19]);
      $fwrite(o, ", %2d", freeNext_memory[20]);
      $fwrite(o, ", %2d", freeNext_memory[21]);
      $fwrite(o, ", %2d", freeNext_memory[22]);
      $fwrite(o, ", %2d", freeNext_memory[23]);
      $fwrite(o, ", %2d", freeNext_memory[24]);
      $fwrite(o, ", %2d", freeNext_memory[25]);
      $fwrite(o, ", %2d", freeNext_memory[26]);
      $fwrite(o, ", %2d", freeNext_memory[27]);
      $fwrite(o, ", %2d", freeNext_memory[28]);
      $fwrite(o, ", %2d", freeNext_memory[29]);
      $fwrite(o, ", %2d", freeNext_memory[30]);
      $fwrite(o, ", %2d", freeNext_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "freeNext_9", freeNext_9_requestedAt, freeNext_9_finishedAt, freeNext_freeNext_9_returnCode, (freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step), (freeNext_9_requestedAt < freeNext_9_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_freeNext_9_index_194", put_freeNext_9_index_194);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "freeNext_10", freeNext_10_requestedAt, freeNext_10_finishedAt, freeNext_freeNext_10_returnCode, (freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step), (freeNext_10_requestedAt < freeNext_10_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_freeNext_10_index_195", put_freeNext_10_index_195);

      $fwrite(o, "            %-38s = %1d\n", "put_freeNext_10_value_196", put_freeNext_10_value_196);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 3, "stuckSize", 1, stuckSize_pc, stuckSize_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 3, 1);
      $fwrite(o, "        %2d", stuckSize_memory[0]);
      $fwrite(o, ", %2d", stuckSize_memory[1]);
      $fwrite(o, ", %2d", stuckSize_memory[2]);
      $fwrite(o, ", %2d", stuckSize_memory[3]);
      $fwrite(o, ", %2d", stuckSize_memory[4]);
      $fwrite(o, ", %2d", stuckSize_memory[5]);
      $fwrite(o, ", %2d", stuckSize_memory[6]);
      $fwrite(o, ", %2d", stuckSize_memory[7]);
      $fwrite(o, ", %2d", stuckSize_memory[8]);
      $fwrite(o, ", %2d", stuckSize_memory[9]);
      $fwrite(o, ", %2d", stuckSize_memory[10]);
      $fwrite(o, ", %2d", stuckSize_memory[11]);
      $fwrite(o, ", %2d", stuckSize_memory[12]);
      $fwrite(o, ", %2d", stuckSize_memory[13]);
      $fwrite(o, ", %2d", stuckSize_memory[14]);
      $fwrite(o, ", %2d", stuckSize_memory[15]);
      $fwrite(o, ", %2d", stuckSize_memory[16]);
      $fwrite(o, ", %2d", stuckSize_memory[17]);
      $fwrite(o, ", %2d", stuckSize_memory[18]);
      $fwrite(o, ", %2d", stuckSize_memory[19]);
      $fwrite(o, ", %2d", stuckSize_memory[20]);
      $fwrite(o, ", %2d", stuckSize_memory[21]);
      $fwrite(o, ", %2d", stuckSize_memory[22]);
      $fwrite(o, ", %2d", stuckSize_memory[23]);
      $fwrite(o, ", %2d", stuckSize_memory[24]);
      $fwrite(o, ", %2d", stuckSize_memory[25]);
      $fwrite(o, ", %2d", stuckSize_memory[26]);
      $fwrite(o, ", %2d", stuckSize_memory[27]);
      $fwrite(o, ", %2d", stuckSize_memory[28]);
      $fwrite(o, ", %2d", stuckSize_memory[29]);
      $fwrite(o, ", %2d", stuckSize_memory[30]);
      $fwrite(o, ", %2d", stuckSize_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckSize_5", stuckSize_5_requestedAt, stuckSize_5_finishedAt, stuckSize_stuckSize_5_returnCode, (stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step), (stuckSize_5_requestedAt < stuckSize_5_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckSize_5_index_36", put_stuckSize_5_index_36);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckSize_6", stuckSize_6_requestedAt, stuckSize_6_finishedAt, stuckSize_stuckSize_6_returnCode, (stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step), (stuckSize_6_requestedAt < stuckSize_6_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckSize_6_index_37", put_stuckSize_6_index_37);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckSize_6_value_38", put_stuckSize_6_value_38);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 4, "stuckKeys", 1, stuckKeys_pc, stuckKeys_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckKeys_memory[0]);
      $fwrite(o, ", %2d", stuckKeys_memory[1]);
      $fwrite(o, ", %2d", stuckKeys_memory[2]);
      $fwrite(o, ", %2d", stuckKeys_memory[3]);
      $fwrite(o, ", %2d", stuckKeys_memory[4]);
      $fwrite(o, ", %2d", stuckKeys_memory[5]);
      $fwrite(o, ", %2d", stuckKeys_memory[6]);
      $fwrite(o, ", %2d", stuckKeys_memory[7]);
      $fwrite(o, ", %2d", stuckKeys_memory[8]);
      $fwrite(o, ", %2d", stuckKeys_memory[9]);
      $fwrite(o, ", %2d", stuckKeys_memory[10]);
      $fwrite(o, ", %2d", stuckKeys_memory[11]);
      $fwrite(o, ", %2d", stuckKeys_memory[12]);
      $fwrite(o, ", %2d", stuckKeys_memory[13]);
      $fwrite(o, ", %2d", stuckKeys_memory[14]);
      $fwrite(o, ", %2d", stuckKeys_memory[15]);
      $fwrite(o, ", %2d", stuckKeys_memory[16]);
      $fwrite(o, ", %2d", stuckKeys_memory[17]);
      $fwrite(o, ", %2d", stuckKeys_memory[18]);
      $fwrite(o, ", %2d", stuckKeys_memory[19]);
      $fwrite(o, ", %2d", stuckKeys_memory[20]);
      $fwrite(o, ", %2d", stuckKeys_memory[21]);
      $fwrite(o, ", %2d", stuckKeys_memory[22]);
      $fwrite(o, ", %2d", stuckKeys_memory[23]);
      $fwrite(o, ", %2d", stuckKeys_memory[24]);
      $fwrite(o, ", %2d", stuckKeys_memory[25]);
      $fwrite(o, ", %2d", stuckKeys_memory[26]);
      $fwrite(o, ", %2d", stuckKeys_memory[27]);
      $fwrite(o, ", %2d", stuckKeys_memory[28]);
      $fwrite(o, ", %2d", stuckKeys_memory[29]);
      $fwrite(o, ", %2d", stuckKeys_memory[30]);
      $fwrite(o, ", %2d", stuckKeys_memory[31]);
      $fwrite(o, ", %2d", stuckKeys_memory[32]);
      $fwrite(o, ", %2d", stuckKeys_memory[33]);
      $fwrite(o, ", %2d", stuckKeys_memory[34]);
      $fwrite(o, ", %2d", stuckKeys_memory[35]);
      $fwrite(o, ", %2d", stuckKeys_memory[36]);
      $fwrite(o, ", %2d", stuckKeys_memory[37]);
      $fwrite(o, ", %2d", stuckKeys_memory[38]);
      $fwrite(o, ", %2d", stuckKeys_memory[39]);
      $fwrite(o, ", %2d", stuckKeys_memory[40]);
      $fwrite(o, ", %2d", stuckKeys_memory[41]);
      $fwrite(o, ", %2d", stuckKeys_memory[42]);
      $fwrite(o, ", %2d", stuckKeys_memory[43]);
      $fwrite(o, ", %2d", stuckKeys_memory[44]);
      $fwrite(o, ", %2d", stuckKeys_memory[45]);
      $fwrite(o, ", %2d", stuckKeys_memory[46]);
      $fwrite(o, ", %2d", stuckKeys_memory[47]);
      $fwrite(o, ", %2d", stuckKeys_memory[48]);
      $fwrite(o, ", %2d", stuckKeys_memory[49]);
      $fwrite(o, ", %2d", stuckKeys_memory[50]);
      $fwrite(o, ", %2d", stuckKeys_memory[51]);
      $fwrite(o, ", %2d", stuckKeys_memory[52]);
      $fwrite(o, ", %2d", stuckKeys_memory[53]);
      $fwrite(o, ", %2d", stuckKeys_memory[54]);
      $fwrite(o, ", %2d", stuckKeys_memory[55]);
      $fwrite(o, ", %2d", stuckKeys_memory[56]);
      $fwrite(o, ", %2d", stuckKeys_memory[57]);
      $fwrite(o, ", %2d", stuckKeys_memory[58]);
      $fwrite(o, ", %2d", stuckKeys_memory[59]);
      $fwrite(o, ", %2d", stuckKeys_memory[60]);
      $fwrite(o, ", %2d", stuckKeys_memory[61]);
      $fwrite(o, ", %2d", stuckKeys_memory[62]);
      $fwrite(o, ", %2d", stuckKeys_memory[63]);
      $fwrite(o, ", %2d", stuckKeys_memory[64]);
      $fwrite(o, ", %2d", stuckKeys_memory[65]);
      $fwrite(o, ", %2d", stuckKeys_memory[66]);
      $fwrite(o, ", %2d", stuckKeys_memory[67]);
      $fwrite(o, ", %2d", stuckKeys_memory[68]);
      $fwrite(o, ", %2d", stuckKeys_memory[69]);
      $fwrite(o, ", %2d", stuckKeys_memory[70]);
      $fwrite(o, ", %2d", stuckKeys_memory[71]);
      $fwrite(o, ", %2d", stuckKeys_memory[72]);
      $fwrite(o, ", %2d", stuckKeys_memory[73]);
      $fwrite(o, ", %2d", stuckKeys_memory[74]);
      $fwrite(o, ", %2d", stuckKeys_memory[75]);
      $fwrite(o, ", %2d", stuckKeys_memory[76]);
      $fwrite(o, ", %2d", stuckKeys_memory[77]);
      $fwrite(o, ", %2d", stuckKeys_memory[78]);
      $fwrite(o, ", %2d", stuckKeys_memory[79]);
      $fwrite(o, ", %2d", stuckKeys_memory[80]);
      $fwrite(o, ", %2d", stuckKeys_memory[81]);
      $fwrite(o, ", %2d", stuckKeys_memory[82]);
      $fwrite(o, ", %2d", stuckKeys_memory[83]);
      $fwrite(o, ", %2d", stuckKeys_memory[84]);
      $fwrite(o, ", %2d", stuckKeys_memory[85]);
      $fwrite(o, ", %2d", stuckKeys_memory[86]);
      $fwrite(o, ", %2d", stuckKeys_memory[87]);
      $fwrite(o, ", %2d", stuckKeys_memory[88]);
      $fwrite(o, ", %2d", stuckKeys_memory[89]);
      $fwrite(o, ", %2d", stuckKeys_memory[90]);
      $fwrite(o, ", %2d", stuckKeys_memory[91]);
      $fwrite(o, ", %2d", stuckKeys_memory[92]);
      $fwrite(o, ", %2d", stuckKeys_memory[93]);
      $fwrite(o, ", %2d", stuckKeys_memory[94]);
      $fwrite(o, ", %2d", stuckKeys_memory[95]);
      $fwrite(o, ", %2d", stuckKeys_memory[96]);
      $fwrite(o, ", %2d", stuckKeys_memory[97]);
      $fwrite(o, ", %2d", stuckKeys_memory[98]);
      $fwrite(o, ", %2d", stuckKeys_memory[99]);
      $fwrite(o, ", %2d", stuckKeys_memory[100]);
      $fwrite(o, ", %2d", stuckKeys_memory[101]);
      $fwrite(o, ", %2d", stuckKeys_memory[102]);
      $fwrite(o, ", %2d", stuckKeys_memory[103]);
      $fwrite(o, ", %2d", stuckKeys_memory[104]);
      $fwrite(o, ", %2d", stuckKeys_memory[105]);
      $fwrite(o, ", %2d", stuckKeys_memory[106]);
      $fwrite(o, ", %2d", stuckKeys_memory[107]);
      $fwrite(o, ", %2d", stuckKeys_memory[108]);
      $fwrite(o, ", %2d", stuckKeys_memory[109]);
      $fwrite(o, ", %2d", stuckKeys_memory[110]);
      $fwrite(o, ", %2d", stuckKeys_memory[111]);
      $fwrite(o, ", %2d", stuckKeys_memory[112]);
      $fwrite(o, ", %2d", stuckKeys_memory[113]);
      $fwrite(o, ", %2d", stuckKeys_memory[114]);
      $fwrite(o, ", %2d", stuckKeys_memory[115]);
      $fwrite(o, ", %2d", stuckKeys_memory[116]);
      $fwrite(o, ", %2d", stuckKeys_memory[117]);
      $fwrite(o, ", %2d", stuckKeys_memory[118]);
      $fwrite(o, ", %2d", stuckKeys_memory[119]);
      $fwrite(o, ", %2d", stuckKeys_memory[120]);
      $fwrite(o, ", %2d", stuckKeys_memory[121]);
      $fwrite(o, ", %2d", stuckKeys_memory[122]);
      $fwrite(o, ", %2d", stuckKeys_memory[123]);
      $fwrite(o, ", %2d", stuckKeys_memory[124]);
      $fwrite(o, ", %2d", stuckKeys_memory[125]);
      $fwrite(o, ", %2d", stuckKeys_memory[126]);
      $fwrite(o, ", %2d", stuckKeys_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckKeys_1", stuckKeys_1_requestedAt, stuckKeys_1_finishedAt, stuckKeys_stuckKeys_1_returnCode, (stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step), (stuckKeys_1_requestedAt < stuckKeys_1_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_1_index_24", put_stuckKeys_1_index_24);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckKeys_2", stuckKeys_2_requestedAt, stuckKeys_2_finishedAt, stuckKeys_stuckKeys_2_returnCode, (stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step), (stuckKeys_2_requestedAt < stuckKeys_2_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_index_25", put_stuckKeys_2_index_25);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_26", put_stuckKeys_2_value_26);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_27", put_stuckKeys_2_value_27);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_28", put_stuckKeys_2_value_28);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_29", put_stuckKeys_2_value_29);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 5, "stuckData", 1, stuckData_pc, stuckData_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckData_memory[0]);
      $fwrite(o, ", %2d", stuckData_memory[1]);
      $fwrite(o, ", %2d", stuckData_memory[2]);
      $fwrite(o, ", %2d", stuckData_memory[3]);
      $fwrite(o, ", %2d", stuckData_memory[4]);
      $fwrite(o, ", %2d", stuckData_memory[5]);
      $fwrite(o, ", %2d", stuckData_memory[6]);
      $fwrite(o, ", %2d", stuckData_memory[7]);
      $fwrite(o, ", %2d", stuckData_memory[8]);
      $fwrite(o, ", %2d", stuckData_memory[9]);
      $fwrite(o, ", %2d", stuckData_memory[10]);
      $fwrite(o, ", %2d", stuckData_memory[11]);
      $fwrite(o, ", %2d", stuckData_memory[12]);
      $fwrite(o, ", %2d", stuckData_memory[13]);
      $fwrite(o, ", %2d", stuckData_memory[14]);
      $fwrite(o, ", %2d", stuckData_memory[15]);
      $fwrite(o, ", %2d", stuckData_memory[16]);
      $fwrite(o, ", %2d", stuckData_memory[17]);
      $fwrite(o, ", %2d", stuckData_memory[18]);
      $fwrite(o, ", %2d", stuckData_memory[19]);
      $fwrite(o, ", %2d", stuckData_memory[20]);
      $fwrite(o, ", %2d", stuckData_memory[21]);
      $fwrite(o, ", %2d", stuckData_memory[22]);
      $fwrite(o, ", %2d", stuckData_memory[23]);
      $fwrite(o, ", %2d", stuckData_memory[24]);
      $fwrite(o, ", %2d", stuckData_memory[25]);
      $fwrite(o, ", %2d", stuckData_memory[26]);
      $fwrite(o, ", %2d", stuckData_memory[27]);
      $fwrite(o, ", %2d", stuckData_memory[28]);
      $fwrite(o, ", %2d", stuckData_memory[29]);
      $fwrite(o, ", %2d", stuckData_memory[30]);
      $fwrite(o, ", %2d", stuckData_memory[31]);
      $fwrite(o, ", %2d", stuckData_memory[32]);
      $fwrite(o, ", %2d", stuckData_memory[33]);
      $fwrite(o, ", %2d", stuckData_memory[34]);
      $fwrite(o, ", %2d", stuckData_memory[35]);
      $fwrite(o, ", %2d", stuckData_memory[36]);
      $fwrite(o, ", %2d", stuckData_memory[37]);
      $fwrite(o, ", %2d", stuckData_memory[38]);
      $fwrite(o, ", %2d", stuckData_memory[39]);
      $fwrite(o, ", %2d", stuckData_memory[40]);
      $fwrite(o, ", %2d", stuckData_memory[41]);
      $fwrite(o, ", %2d", stuckData_memory[42]);
      $fwrite(o, ", %2d", stuckData_memory[43]);
      $fwrite(o, ", %2d", stuckData_memory[44]);
      $fwrite(o, ", %2d", stuckData_memory[45]);
      $fwrite(o, ", %2d", stuckData_memory[46]);
      $fwrite(o, ", %2d", stuckData_memory[47]);
      $fwrite(o, ", %2d", stuckData_memory[48]);
      $fwrite(o, ", %2d", stuckData_memory[49]);
      $fwrite(o, ", %2d", stuckData_memory[50]);
      $fwrite(o, ", %2d", stuckData_memory[51]);
      $fwrite(o, ", %2d", stuckData_memory[52]);
      $fwrite(o, ", %2d", stuckData_memory[53]);
      $fwrite(o, ", %2d", stuckData_memory[54]);
      $fwrite(o, ", %2d", stuckData_memory[55]);
      $fwrite(o, ", %2d", stuckData_memory[56]);
      $fwrite(o, ", %2d", stuckData_memory[57]);
      $fwrite(o, ", %2d", stuckData_memory[58]);
      $fwrite(o, ", %2d", stuckData_memory[59]);
      $fwrite(o, ", %2d", stuckData_memory[60]);
      $fwrite(o, ", %2d", stuckData_memory[61]);
      $fwrite(o, ", %2d", stuckData_memory[62]);
      $fwrite(o, ", %2d", stuckData_memory[63]);
      $fwrite(o, ", %2d", stuckData_memory[64]);
      $fwrite(o, ", %2d", stuckData_memory[65]);
      $fwrite(o, ", %2d", stuckData_memory[66]);
      $fwrite(o, ", %2d", stuckData_memory[67]);
      $fwrite(o, ", %2d", stuckData_memory[68]);
      $fwrite(o, ", %2d", stuckData_memory[69]);
      $fwrite(o, ", %2d", stuckData_memory[70]);
      $fwrite(o, ", %2d", stuckData_memory[71]);
      $fwrite(o, ", %2d", stuckData_memory[72]);
      $fwrite(o, ", %2d", stuckData_memory[73]);
      $fwrite(o, ", %2d", stuckData_memory[74]);
      $fwrite(o, ", %2d", stuckData_memory[75]);
      $fwrite(o, ", %2d", stuckData_memory[76]);
      $fwrite(o, ", %2d", stuckData_memory[77]);
      $fwrite(o, ", %2d", stuckData_memory[78]);
      $fwrite(o, ", %2d", stuckData_memory[79]);
      $fwrite(o, ", %2d", stuckData_memory[80]);
      $fwrite(o, ", %2d", stuckData_memory[81]);
      $fwrite(o, ", %2d", stuckData_memory[82]);
      $fwrite(o, ", %2d", stuckData_memory[83]);
      $fwrite(o, ", %2d", stuckData_memory[84]);
      $fwrite(o, ", %2d", stuckData_memory[85]);
      $fwrite(o, ", %2d", stuckData_memory[86]);
      $fwrite(o, ", %2d", stuckData_memory[87]);
      $fwrite(o, ", %2d", stuckData_memory[88]);
      $fwrite(o, ", %2d", stuckData_memory[89]);
      $fwrite(o, ", %2d", stuckData_memory[90]);
      $fwrite(o, ", %2d", stuckData_memory[91]);
      $fwrite(o, ", %2d", stuckData_memory[92]);
      $fwrite(o, ", %2d", stuckData_memory[93]);
      $fwrite(o, ", %2d", stuckData_memory[94]);
      $fwrite(o, ", %2d", stuckData_memory[95]);
      $fwrite(o, ", %2d", stuckData_memory[96]);
      $fwrite(o, ", %2d", stuckData_memory[97]);
      $fwrite(o, ", %2d", stuckData_memory[98]);
      $fwrite(o, ", %2d", stuckData_memory[99]);
      $fwrite(o, ", %2d", stuckData_memory[100]);
      $fwrite(o, ", %2d", stuckData_memory[101]);
      $fwrite(o, ", %2d", stuckData_memory[102]);
      $fwrite(o, ", %2d", stuckData_memory[103]);
      $fwrite(o, ", %2d", stuckData_memory[104]);
      $fwrite(o, ", %2d", stuckData_memory[105]);
      $fwrite(o, ", %2d", stuckData_memory[106]);
      $fwrite(o, ", %2d", stuckData_memory[107]);
      $fwrite(o, ", %2d", stuckData_memory[108]);
      $fwrite(o, ", %2d", stuckData_memory[109]);
      $fwrite(o, ", %2d", stuckData_memory[110]);
      $fwrite(o, ", %2d", stuckData_memory[111]);
      $fwrite(o, ", %2d", stuckData_memory[112]);
      $fwrite(o, ", %2d", stuckData_memory[113]);
      $fwrite(o, ", %2d", stuckData_memory[114]);
      $fwrite(o, ", %2d", stuckData_memory[115]);
      $fwrite(o, ", %2d", stuckData_memory[116]);
      $fwrite(o, ", %2d", stuckData_memory[117]);
      $fwrite(o, ", %2d", stuckData_memory[118]);
      $fwrite(o, ", %2d", stuckData_memory[119]);
      $fwrite(o, ", %2d", stuckData_memory[120]);
      $fwrite(o, ", %2d", stuckData_memory[121]);
      $fwrite(o, ", %2d", stuckData_memory[122]);
      $fwrite(o, ", %2d", stuckData_memory[123]);
      $fwrite(o, ", %2d", stuckData_memory[124]);
      $fwrite(o, ", %2d", stuckData_memory[125]);
      $fwrite(o, ", %2d", stuckData_memory[126]);
      $fwrite(o, ", %2d", stuckData_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckData_3", stuckData_3_requestedAt, stuckData_3_finishedAt, stuckData_stuckData_3_returnCode, (stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step), (stuckData_3_requestedAt < stuckData_3_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_3_index_30", put_stuckData_3_index_30);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckData_4", stuckData_4_requestedAt, stuckData_4_finishedAt, stuckData_stuckData_4_returnCode, (stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step), (stuckData_4_requestedAt < stuckData_4_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_index_31", put_stuckData_4_index_31);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_32", put_stuckData_4_value_32);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_33", put_stuckData_4_value_33);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_34", put_stuckData_4_value_34);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_35", put_stuckData_4_value_35);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 6, "put", 984, put_pc, put_returnCode);
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_k_0", put_k_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_d_1", put_d_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_2", put_i_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_l_3", put_l_3);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_4", put_index_4);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_5", put_size_5);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_6", put_isLeaf_6);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_7", put_nextFree_7);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_8", put_Key_0_8);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_9", put_KeyCompares_0_9);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_10", put_KeyCollapse_0_10);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_11", put_Data_0_11);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_12", put_Key_1_12);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_13", put_KeyCompares_1_13);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_14", put_KeyCollapse_1_14);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_15", put_Data_1_15);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_16", put_Key_2_16);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_17", put_KeyCompares_2_17);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_18", put_KeyCollapse_2_18);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_19", put_Data_2_19);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_20", put_Key_3_20);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_21", put_KeyCompares_3_21);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_22", put_KeyCollapse_3_22);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_23", put_Data_3_23);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_1_index_24", put_stuckKeys_1_index_24);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_index_25", put_stuckKeys_2_index_25);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_26", put_stuckKeys_2_value_26);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_27", put_stuckKeys_2_value_27);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_28", put_stuckKeys_2_value_28);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_29", put_stuckKeys_2_value_29);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_3_index_30", put_stuckData_3_index_30);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_index_31", put_stuckData_4_index_31);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_32", put_stuckData_4_value_32);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_33", put_stuckData_4_value_33);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_34", put_stuckData_4_value_34);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_35", put_stuckData_4_value_35);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckSize_5_index_36", put_stuckSize_5_index_36);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckSize_6_index_37", put_stuckSize_6_index_37);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckSize_6_value_38", put_stuckSize_6_value_38);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsLeaf_7_index_39", put_stuckIsLeaf_7_index_39);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsLeaf_8_index_40", put_stuckIsLeaf_8_index_40);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsLeaf_8_value_41", put_stuckIsLeaf_8_value_41);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_42", put_Found_42);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_43", put_Key_43);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_44", put_FoundKey_44);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_45", put_Data_45);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_46", put_BtreeIndex_46);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_47", put_StuckIndex_47);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_48", put_MergeSuccess_48);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_49", put_index_49);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_50", put_size_50);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_51", put_isLeaf_51);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_52", put_nextFree_52);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_53", put_Key_0_53);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_54", put_KeyCompares_0_54);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_55", put_KeyCollapse_0_55);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_56", put_Data_0_56);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_57", put_Key_1_57);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_58", put_KeyCompares_1_58);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_59", put_KeyCollapse_1_59);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_60", put_Data_1_60);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_61", put_Key_2_61);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_62", put_KeyCompares_2_62);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_63", put_KeyCollapse_2_63);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_64", put_Data_2_64);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_65", put_Key_3_65);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_66", put_KeyCompares_3_66);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_67", put_KeyCollapse_3_67);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_68", put_Data_3_68);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_69", put_Found_69);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_70", put_Key_70);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_71", put_FoundKey_71);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_72", put_Data_72);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_73", put_BtreeIndex_73);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_74", put_StuckIndex_74);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_75", put_MergeSuccess_75);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_76", put_index_76);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_77", put_size_77);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_78", put_isLeaf_78);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_79", put_nextFree_79);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_80", put_Key_0_80);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_81", put_KeyCompares_0_81);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_82", put_KeyCollapse_0_82);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_83", put_Data_0_83);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_84", put_Key_1_84);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_85", put_KeyCompares_1_85);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_86", put_KeyCollapse_1_86);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_87", put_Data_1_87);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_88", put_Key_2_88);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_89", put_KeyCompares_2_89);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_90", put_KeyCollapse_2_90);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_91", put_Data_2_91);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_92", put_Key_3_92);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_93", put_KeyCompares_3_93);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_94", put_KeyCollapse_3_94);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_95", put_Data_3_95);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_96", put_Found_96);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_97", put_Key_97);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_98", put_FoundKey_98);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_99", put_Data_99);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_100", put_BtreeIndex_100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_101", put_StuckIndex_101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_102", put_MergeSuccess_102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_child_103", put_child_103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_parent_104", put_parent_104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childInparent_105", put_childInparent_105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_found_106", put_found_106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_full_107", put_full_107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_108", put_i_108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_notFull_109", put_notFull_109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_110", put_index_110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_111", put_size_111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_112", put_isLeaf_112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_113", put_nextFree_113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_114", put_Key_0_114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_115", put_KeyCompares_0_115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_116", put_KeyCollapse_0_116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_117", put_Data_0_117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_118", put_Key_1_118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_119", put_KeyCompares_1_119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_120", put_KeyCollapse_1_120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_121", put_Data_1_121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_122", put_Key_2_122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_123", put_KeyCompares_2_123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_124", put_KeyCollapse_2_124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_125", put_Data_2_125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_126", put_Key_3_126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_127", put_KeyCompares_3_127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_128", put_KeyCollapse_3_128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_129", put_Data_3_129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_130", put_Found_130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_131", put_Key_131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_132", put_FoundKey_132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_133", put_Data_133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_134", put_BtreeIndex_134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_135", put_StuckIndex_135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_136", put_MergeSuccess_136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_137", put_index_137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_138", put_size_138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_139", put_isLeaf_139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_140", put_nextFree_140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_141", put_Key_0_141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_142", put_KeyCompares_0_142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_143", put_KeyCollapse_0_143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_144", put_Data_0_144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_145", put_Key_1_145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_146", put_KeyCompares_1_146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_147", put_KeyCollapse_1_147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_148", put_Data_1_148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_149", put_Key_2_149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_150", put_KeyCompares_2_150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_151", put_KeyCollapse_2_151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_152", put_Data_2_152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_153", put_Key_3_153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_154", put_KeyCompares_3_154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_155", put_KeyCollapse_3_155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_156", put_Data_3_156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_157", put_Found_157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_158", put_Key_158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_159", put_FoundKey_159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_160", put_Data_160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_161", put_BtreeIndex_161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_162", put_StuckIndex_162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_163", put_MergeSuccess_163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_164", put_index_164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_165", put_size_165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_166", put_isLeaf_166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_167", put_nextFree_167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_168", put_Key_0_168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_169", put_KeyCompares_0_169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_170", put_KeyCollapse_0_170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_171", put_Data_0_171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_172", put_Key_1_172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_173", put_KeyCompares_1_173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_174", put_KeyCollapse_1_174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_175", put_Data_1_175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_176", put_Key_2_176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_177", put_KeyCompares_2_177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_178", put_KeyCollapse_2_178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_179", put_Data_2_179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_180", put_Key_3_180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_181", put_KeyCompares_3_181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_182", put_KeyCollapse_3_182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_183", put_Data_3_183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_184", put_Found_184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_185", put_Key_185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_186", put_FoundKey_186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_187", put_Data_187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_188", put_BtreeIndex_188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_189", put_StuckIndex_189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_190", put_MergeSuccess_190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_191", put_indexLeft_191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_192", put_indexRight_192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_193", put_midKey_193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_freeNext_9_index_194", put_freeNext_9_index_194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_freeNext_10_index_195", put_freeNext_10_index_195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_freeNext_10_value_196", put_freeNext_10_value_196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsFree_11_index_197", put_stuckIsFree_11_index_197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsFree_11_value_198", put_stuckIsFree_11_value_198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_199", put_root_199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_200", put_next_200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_201", put_isLeaf_201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_202", put_isFree_202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_203", put_root_203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_204", put_next_204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_205", put_isLeaf_205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_206", put_isFree_206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_207", put_i_207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_notFull_208", put_notFull_208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_209", put_index_209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_210", put_size_210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_211", put_isLeaf_211);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_212", put_nextFree_212);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_213", put_Key_0_213);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_214", put_KeyCompares_0_214);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_215", put_KeyCollapse_0_215);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_216", put_Data_0_216);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_217", put_Key_1_217);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_218", put_KeyCompares_1_218);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_219", put_KeyCollapse_1_219);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_220", put_Data_1_220);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_221", put_Key_2_221);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_222", put_KeyCompares_2_222);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_223", put_KeyCollapse_2_223);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_224", put_Data_2_224);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_225", put_Key_3_225);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_226", put_KeyCompares_3_226);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_227", put_KeyCollapse_3_227);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_228", put_Data_3_228);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_229", put_Found_229);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_230", put_Key_230);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_231", put_FoundKey_231);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_232", put_Data_232);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_233", put_BtreeIndex_233);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_234", put_StuckIndex_234);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_235", put_MergeSuccess_235);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_236", put_index_236);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_237", put_size_237);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_238", put_isLeaf_238);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_239", put_nextFree_239);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_240", put_Key_0_240);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_241", put_KeyCompares_0_241);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_242", put_KeyCollapse_0_242);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_243", put_Data_0_243);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_244", put_Key_1_244);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_245", put_KeyCompares_1_245);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_246", put_KeyCollapse_1_246);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_247", put_Data_1_247);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_248", put_Key_2_248);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_249", put_KeyCompares_2_249);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_250", put_KeyCollapse_2_250);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_251", put_Data_2_251);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_252", put_Key_3_252);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_253", put_KeyCompares_3_253);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_254", put_KeyCollapse_3_254);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_255", put_Data_3_255);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_256", put_Found_256);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_257", put_Key_257);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_258", put_FoundKey_258);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_259", put_Data_259);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_260", put_BtreeIndex_260);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_261", put_StuckIndex_261);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_262", put_MergeSuccess_262);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_263", put_index_263);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_264", put_size_264);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_265", put_isLeaf_265);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_266", put_nextFree_266);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_267", put_Key_0_267);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_268", put_KeyCompares_0_268);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_269", put_KeyCollapse_0_269);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_270", put_Data_0_270);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_271", put_Key_1_271);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_272", put_KeyCompares_1_272);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_273", put_KeyCollapse_1_273);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_274", put_Data_1_274);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_275", put_Key_2_275);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_276", put_KeyCompares_2_276);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_277", put_KeyCollapse_2_277);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_278", put_Data_2_278);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_279", put_Key_3_279);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_280", put_KeyCompares_3_280);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_281", put_KeyCollapse_3_281);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_282", put_Data_3_282);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_283", put_Found_283);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_284", put_Key_284);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_285", put_FoundKey_285);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_286", put_Data_286);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_287", put_BtreeIndex_287);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_288", put_StuckIndex_288);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_289", put_MergeSuccess_289);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_290", put_indexLeft_290);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_291", put_indexRight_291);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_292", put_midKey_292);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_293", put_root_293);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_294", put_next_294);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_295", put_isLeaf_295);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_296", put_isFree_296);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_297", put_root_297);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_298", put_next_298);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_299", put_isLeaf_299);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_300", put_isFree_300);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_301", put_index_301);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_302", put_size_302);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_303", put_isLeaf_303);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_304", put_nextFree_304);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_305", put_Key_0_305);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_306", put_KeyCompares_0_306);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_307", put_KeyCollapse_0_307);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_308", put_Data_0_308);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_309", put_Key_1_309);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_310", put_KeyCompares_1_310);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_311", put_KeyCollapse_1_311);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_312", put_Data_1_312);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_313", put_Key_2_313);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_314", put_KeyCompares_2_314);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_315", put_KeyCollapse_2_315);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_316", put_Data_2_316);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_317", put_Key_3_317);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_318", put_KeyCompares_3_318);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_319", put_KeyCollapse_3_319);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_320", put_Data_3_320);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_321", put_Found_321);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_322", put_Key_322);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_323", put_FoundKey_323);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_324", put_Data_324);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_325", put_BtreeIndex_325);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_326", put_StuckIndex_326);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_327", put_MergeSuccess_327);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_328", put_index_328);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_329", put_size_329);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_330", put_isLeaf_330);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_331", put_nextFree_331);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_332", put_Key_0_332);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_333", put_KeyCompares_0_333);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_334", put_KeyCollapse_0_334);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_335", put_Data_0_335);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_336", put_Key_1_336);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_337", put_KeyCompares_1_337);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_338", put_KeyCollapse_1_338);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_339", put_Data_1_339);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_340", put_Key_2_340);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_341", put_KeyCompares_2_341);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_342", put_KeyCollapse_2_342);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_343", put_Data_2_343);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_344", put_Key_3_344);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_345", put_KeyCompares_3_345);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_346", put_KeyCollapse_3_346);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_347", put_Data_3_347);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_348", put_Found_348);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_349", put_Key_349);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_350", put_FoundKey_350);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_351", put_Data_351);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_352", put_BtreeIndex_352);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_353", put_StuckIndex_353);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_354", put_MergeSuccess_354);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_355", put_index_355);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_356", put_size_356);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_357", put_isLeaf_357);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_358", put_nextFree_358);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_359", put_Key_0_359);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_360", put_KeyCompares_0_360);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_361", put_KeyCollapse_0_361);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_362", put_Data_0_362);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_363", put_Key_1_363);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_364", put_KeyCompares_1_364);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_365", put_KeyCollapse_1_365);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_366", put_Data_1_366);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_367", put_Key_2_367);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_368", put_KeyCompares_2_368);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_369", put_KeyCollapse_2_369);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_370", put_Data_2_370);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_371", put_Key_3_371);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_372", put_KeyCompares_3_372);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_373", put_KeyCollapse_3_373);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_374", put_Data_3_374);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_375", put_Found_375);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_376", put_Key_376);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_377", put_FoundKey_377);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_378", put_Data_378);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_379", put_BtreeIndex_379);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_380", put_StuckIndex_380);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_381", put_MergeSuccess_381);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_382", put_index_382);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_383", put_size_383);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_384", put_isLeaf_384);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_385", put_nextFree_385);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_386", put_Key_0_386);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_387", put_KeyCompares_0_387);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_388", put_KeyCollapse_0_388);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_389", put_Data_0_389);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_390", put_Key_1_390);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_391", put_KeyCompares_1_391);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_392", put_KeyCollapse_1_392);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_393", put_Data_1_393);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_394", put_Key_2_394);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_395", put_KeyCompares_2_395);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_396", put_KeyCollapse_2_396);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_397", put_Data_2_397);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_398", put_Key_3_398);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_399", put_KeyCompares_3_399);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_400", put_KeyCollapse_3_400);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_401", put_Data_3_401);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_402", put_Found_402);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_403", put_Key_403);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_404", put_FoundKey_404);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_405", put_Data_405);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_406", put_BtreeIndex_406);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_407", put_StuckIndex_407);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_408", put_MergeSuccess_408);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_409", put_childKey_409);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_410", put_childData_410);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_411", put_indexLeft_411);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_412", put_indexRight_412);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_413", put_midKey_413);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_414", put_root_414);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_415", put_next_415);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_416", put_isLeaf_416);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_417", put_isFree_417);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_418", put_index_418);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_419", put_size_419);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_420", put_isLeaf_420);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_421", put_nextFree_421);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_422", put_Key_0_422);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_423", put_KeyCompares_0_423);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_424", put_KeyCollapse_0_424);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_425", put_Data_0_425);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_426", put_Key_1_426);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_427", put_KeyCompares_1_427);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_428", put_KeyCollapse_1_428);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_429", put_Data_1_429);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_430", put_Key_2_430);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_431", put_KeyCompares_2_431);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_432", put_KeyCollapse_2_432);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_433", put_Data_2_433);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_434", put_Key_3_434);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_435", put_KeyCompares_3_435);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_436", put_KeyCollapse_3_436);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_437", put_Data_3_437);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_438", put_Found_438);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_439", put_Key_439);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_440", put_FoundKey_440);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_441", put_Data_441);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_442", put_BtreeIndex_442);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_443", put_StuckIndex_443);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_444", put_MergeSuccess_444);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_445", put_index_445);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_446", put_size_446);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_447", put_isLeaf_447);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_448", put_nextFree_448);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_449", put_Key_0_449);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_450", put_KeyCompares_0_450);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_451", put_KeyCollapse_0_451);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_452", put_Data_0_452);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_453", put_Key_1_453);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_454", put_KeyCompares_1_454);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_455", put_KeyCollapse_1_455);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_456", put_Data_1_456);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_457", put_Key_2_457);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_458", put_KeyCompares_2_458);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_459", put_KeyCollapse_2_459);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_460", put_Data_2_460);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_461", put_Key_3_461);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_462", put_KeyCompares_3_462);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_463", put_KeyCollapse_3_463);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_464", put_Data_3_464);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_465", put_Found_465);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_466", put_Key_466);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_467", put_FoundKey_467);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_468", put_Data_468);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_469", put_BtreeIndex_469);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_470", put_StuckIndex_470);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_471", put_MergeSuccess_471);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_472", put_index_472);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_473", put_size_473);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_474", put_isLeaf_474);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_475", put_nextFree_475);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_476", put_Key_0_476);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_477", put_KeyCompares_0_477);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_478", put_KeyCollapse_0_478);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_479", put_Data_0_479);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_480", put_Key_1_480);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_481", put_KeyCompares_1_481);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_482", put_KeyCollapse_1_482);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_483", put_Data_1_483);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_484", put_Key_2_484);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_485", put_KeyCompares_2_485);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_486", put_KeyCollapse_2_486);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_487", put_Data_2_487);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_488", put_Key_3_488);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_489", put_KeyCompares_3_489);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_490", put_KeyCollapse_3_490);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_491", put_Data_3_491);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_492", put_Found_492);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_493", put_Key_493);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_494", put_FoundKey_494);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_495", put_Data_495);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_496", put_BtreeIndex_496);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_497", put_StuckIndex_497);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_498", put_MergeSuccess_498);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childIndex_499", put_childIndex_499);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_leftIndex_500", put_leftIndex_500);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_501", put_midKey_501);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_502", put_root_502);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_503", put_next_503);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_504", put_isLeaf_504);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_505", put_isFree_505);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_506", put_i_506);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_notFull_507", put_notFull_507);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_508", put_index_508);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_509", put_size_509);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_510", put_isLeaf_510);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_511", put_nextFree_511);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_512", put_Key_0_512);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_513", put_KeyCompares_0_513);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_514", put_KeyCollapse_0_514);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_515", put_Data_0_515);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_516", put_Key_1_516);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_517", put_KeyCompares_1_517);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_518", put_KeyCollapse_1_518);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_519", put_Data_1_519);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_520", put_Key_2_520);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_521", put_KeyCompares_2_521);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_522", put_KeyCollapse_2_522);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_523", put_Data_2_523);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_524", put_Key_3_524);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_525", put_KeyCompares_3_525);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_526", put_KeyCollapse_3_526);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_527", put_Data_3_527);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_528", put_Found_528);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_529", put_Key_529);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_530", put_FoundKey_530);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_531", put_Data_531);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_532", put_BtreeIndex_532);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_533", put_StuckIndex_533);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_534", put_MergeSuccess_534);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_535", put_index_535);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_536", put_size_536);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_537", put_isLeaf_537);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_538", put_nextFree_538);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_539", put_Key_0_539);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_540", put_KeyCompares_0_540);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_541", put_KeyCollapse_0_541);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_542", put_Data_0_542);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_543", put_Key_1_543);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_544", put_KeyCompares_1_544);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_545", put_KeyCollapse_1_545);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_546", put_Data_1_546);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_547", put_Key_2_547);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_548", put_KeyCompares_2_548);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_549", put_KeyCollapse_2_549);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_550", put_Data_2_550);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_551", put_Key_3_551);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_552", put_KeyCompares_3_552);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_553", put_KeyCollapse_3_553);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_554", put_Data_3_554);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_555", put_Found_555);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_556", put_Key_556);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_557", put_FoundKey_557);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_558", put_Data_558);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_559", put_BtreeIndex_559);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_560", put_StuckIndex_560);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_561", put_MergeSuccess_561);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_562", put_index_562);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_563", put_size_563);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_564", put_isLeaf_564);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_565", put_nextFree_565);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_566", put_Key_0_566);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_567", put_KeyCompares_0_567);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_568", put_KeyCollapse_0_568);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_569", put_Data_0_569);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_570", put_Key_1_570);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_571", put_KeyCompares_1_571);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_572", put_KeyCollapse_1_572);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_573", put_Data_1_573);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_574", put_Key_2_574);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_575", put_KeyCompares_2_575);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_576", put_KeyCollapse_2_576);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_577", put_Data_2_577);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_578", put_Key_3_578);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_579", put_KeyCompares_3_579);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_580", put_KeyCollapse_3_580);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_581", put_Data_3_581);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_582", put_Found_582);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_583", put_Key_583);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_584", put_FoundKey_584);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_585", put_Data_585);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_586", put_BtreeIndex_586);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_587", put_StuckIndex_587);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_588", put_MergeSuccess_588);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_589", put_index_589);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_590", put_size_590);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_591", put_isLeaf_591);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_592", put_nextFree_592);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_593", put_Key_0_593);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_594", put_KeyCompares_0_594);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_595", put_KeyCollapse_0_595);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_596", put_Data_0_596);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_597", put_Key_1_597);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_598", put_KeyCompares_1_598);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_599", put_KeyCollapse_1_599);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_600", put_Data_1_600);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_601", put_Key_2_601);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_602", put_KeyCompares_2_602);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_603", put_KeyCollapse_2_603);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_604", put_Data_2_604);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_605", put_Key_3_605);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_606", put_KeyCompares_3_606);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_607", put_KeyCollapse_3_607);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_608", put_Data_3_608);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_609", put_Found_609);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_610", put_Key_610);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_611", put_FoundKey_611);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_612", put_Data_612);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_613", put_BtreeIndex_613);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_614", put_StuckIndex_614);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_615", put_MergeSuccess_615);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_616", put_childKey_616);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_617", put_childData_617);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_618", put_indexLeft_618);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_619", put_indexRight_619);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_620", put_midKey_620);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_621", put_root_621);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_622", put_next_622);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_623", put_isLeaf_623);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_624", put_isFree_624);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_625", put_index_625);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_626", put_size_626);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_627", put_isLeaf_627);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_628", put_nextFree_628);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_629", put_Key_0_629);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_630", put_KeyCompares_0_630);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_631", put_KeyCollapse_0_631);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_632", put_Data_0_632);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_633", put_Key_1_633);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_634", put_KeyCompares_1_634);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_635", put_KeyCollapse_1_635);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_636", put_Data_1_636);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_637", put_Key_2_637);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_638", put_KeyCompares_2_638);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_639", put_KeyCollapse_2_639);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_640", put_Data_2_640);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_641", put_Key_3_641);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_642", put_KeyCompares_3_642);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_643", put_KeyCollapse_3_643);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_644", put_Data_3_644);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_645", put_Found_645);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_646", put_Key_646);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_647", put_FoundKey_647);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_648", put_Data_648);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_649", put_BtreeIndex_649);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_650", put_StuckIndex_650);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_651", put_MergeSuccess_651);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_652", put_index_652);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_653", put_size_653);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_654", put_isLeaf_654);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_655", put_nextFree_655);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_656", put_Key_0_656);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_657", put_KeyCompares_0_657);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_658", put_KeyCollapse_0_658);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_659", put_Data_0_659);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_660", put_Key_1_660);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_661", put_KeyCompares_1_661);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_662", put_KeyCollapse_1_662);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_663", put_Data_1_663);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_664", put_Key_2_664);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_665", put_KeyCompares_2_665);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_666", put_KeyCollapse_2_666);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_667", put_Data_2_667);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_668", put_Key_3_668);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_669", put_KeyCompares_3_669);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_670", put_KeyCollapse_3_670);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_671", put_Data_3_671);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_672", put_Found_672);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_673", put_Key_673);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_674", put_FoundKey_674);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_675", put_Data_675);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_676", put_BtreeIndex_676);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_677", put_StuckIndex_677);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_678", put_MergeSuccess_678);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_679", put_index_679);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_680", put_size_680);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_681", put_isLeaf_681);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_682", put_nextFree_682);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_683", put_Key_0_683);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_684", put_KeyCompares_0_684);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_685", put_KeyCollapse_0_685);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_686", put_Data_0_686);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_687", put_Key_1_687);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_688", put_KeyCompares_1_688);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_689", put_KeyCollapse_1_689);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_690", put_Data_1_690);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_691", put_Key_2_691);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_692", put_KeyCompares_2_692);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_693", put_KeyCollapse_2_693);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_694", put_Data_2_694);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_695", put_Key_3_695);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_696", put_KeyCompares_3_696);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_697", put_KeyCollapse_3_697);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_698", put_Data_3_698);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_699", put_Found_699);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_700", put_Key_700);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_701", put_FoundKey_701);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_702", put_Data_702);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_703", put_BtreeIndex_703);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_704", put_StuckIndex_704);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_705", put_MergeSuccess_705);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_706", put_index_706);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_707", put_size_707);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_708", put_isLeaf_708);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_709", put_nextFree_709);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_710", put_Key_0_710);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_711", put_KeyCompares_0_711);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_712", put_KeyCollapse_0_712);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_713", put_Data_0_713);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_714", put_Key_1_714);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_715", put_KeyCompares_1_715);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_716", put_KeyCollapse_1_716);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_717", put_Data_1_717);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_718", put_Key_2_718);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_719", put_KeyCompares_2_719);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_720", put_KeyCollapse_2_720);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_721", put_Data_2_721);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_722", put_Key_3_722);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_723", put_KeyCompares_3_723);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_724", put_KeyCollapse_3_724);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_725", put_Data_3_725);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_726", put_Found_726);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_727", put_Key_727);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_728", put_FoundKey_728);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_729", put_Data_729);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_730", put_BtreeIndex_730);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_731", put_StuckIndex_731);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_732", put_MergeSuccess_732);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_733", put_childKey_733);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_734", put_childData_734);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_735", put_indexLeft_735);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_736", put_indexRight_736);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_737", put_midKey_737);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_738", put_root_738);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_739", put_next_739);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_740", put_isLeaf_740);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_741", put_isFree_741);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_742", put_index_742);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_743", put_size_743);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_744", put_isLeaf_744);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_745", put_nextFree_745);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_746", put_Key_0_746);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_747", put_KeyCompares_0_747);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_748", put_KeyCollapse_0_748);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_749", put_Data_0_749);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_750", put_Key_1_750);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_751", put_KeyCompares_1_751);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_752", put_KeyCollapse_1_752);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_753", put_Data_1_753);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_754", put_Key_2_754);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_755", put_KeyCompares_2_755);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_756", put_KeyCollapse_2_756);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_757", put_Data_2_757);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_758", put_Key_3_758);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_759", put_KeyCompares_3_759);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_760", put_KeyCollapse_3_760);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_761", put_Data_3_761);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_762", put_Found_762);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_763", put_Key_763);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_764", put_FoundKey_764);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_765", put_Data_765);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_766", put_BtreeIndex_766);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_767", put_StuckIndex_767);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_768", put_MergeSuccess_768);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_position_769", put_position_769);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_770", put_index_770);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index1_771", put_index1_771);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_within_772", put_within_772);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_773", put_isLeaf_773);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_774", put_index_774);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_775", put_size_775);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_776", put_isLeaf_776);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_777", put_nextFree_777);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_778", put_Key_0_778);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_779", put_KeyCompares_0_779);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_780", put_KeyCollapse_0_780);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_781", put_Data_0_781);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_782", put_Key_1_782);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_783", put_KeyCompares_1_783);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_784", put_KeyCollapse_1_784);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_785", put_Data_1_785);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_786", put_Key_2_786);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_787", put_KeyCompares_2_787);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_788", put_KeyCollapse_2_788);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_789", put_Data_2_789);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_790", put_Key_3_790);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_791", put_KeyCompares_3_791);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_792", put_KeyCollapse_3_792);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_793", put_Data_3_793);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_794", put_Found_794);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_795", put_Key_795);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_796", put_FoundKey_796);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_797", put_Data_797);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_798", put_BtreeIndex_798);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_799", put_StuckIndex_799);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_800", put_MergeSuccess_800);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_801", put_index_801);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_802", put_size_802);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_803", put_isLeaf_803);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_804", put_nextFree_804);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_805", put_Key_0_805);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_806", put_KeyCompares_0_806);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_807", put_KeyCollapse_0_807);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_808", put_Data_0_808);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_809", put_Key_1_809);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_810", put_KeyCompares_1_810);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_811", put_KeyCollapse_1_811);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_812", put_Data_1_812);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_813", put_Key_2_813);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_814", put_KeyCompares_2_814);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_815", put_KeyCollapse_2_815);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_816", put_Data_2_816);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_817", put_Key_3_817);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_818", put_KeyCompares_3_818);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_819", put_KeyCollapse_3_819);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_820", put_Data_3_820);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_821", put_Found_821);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_822", put_Key_822);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_823", put_FoundKey_823);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_824", put_Data_824);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_825", put_BtreeIndex_825);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_826", put_StuckIndex_826);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_827", put_MergeSuccess_827);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_828", put_index_828);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_829", put_size_829);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_830", put_isLeaf_830);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_831", put_nextFree_831);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_832", put_Key_0_832);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_833", put_KeyCompares_0_833);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_834", put_KeyCollapse_0_834);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_835", put_Data_0_835);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_836", put_Key_1_836);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_837", put_KeyCompares_1_837);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_838", put_KeyCollapse_1_838);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_839", put_Data_1_839);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_840", put_Key_2_840);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_841", put_KeyCompares_2_841);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_842", put_KeyCollapse_2_842);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_843", put_Data_2_843);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_844", put_Key_3_844);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_845", put_KeyCompares_3_845);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_846", put_KeyCollapse_3_846);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_847", put_Data_3_847);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_848", put_Found_848);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_849", put_Key_849);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_850", put_FoundKey_850);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_851", put_Data_851);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_852", put_BtreeIndex_852);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_853", put_StuckIndex_853);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_854", put_MergeSuccess_854);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_855", put_childKey_855);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_856", put_childData_856);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_857", put_indexLeft_857);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_858", put_indexRight_858);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_859", put_midKey_859);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_860", put_success_860);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_861", put_test_861);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_862", put_next_862);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_863", put_root_863);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_864", put_isFree_864);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_865", put_next_865);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_866", put_root_866);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_867", put_isFree_867);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_868", put_index_868);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_869", put_size_869);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_870", put_isLeaf_870);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_871", put_nextFree_871);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_872", put_Key_0_872);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_873", put_KeyCompares_0_873);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_874", put_KeyCollapse_0_874);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_875", put_Data_0_875);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_876", put_Key_1_876);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_877", put_KeyCompares_1_877);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_878", put_KeyCollapse_1_878);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_879", put_Data_1_879);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_880", put_Key_2_880);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_881", put_KeyCompares_2_881);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_882", put_KeyCollapse_2_882);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_883", put_Data_2_883);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_884", put_Key_3_884);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_885", put_KeyCompares_3_885);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_886", put_KeyCollapse_3_886);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_887", put_Data_3_887);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_888", put_Found_888);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_889", put_Key_889);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_890", put_FoundKey_890);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_891", put_Data_891);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_892", put_BtreeIndex_892);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_893", put_StuckIndex_893);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_894", put_MergeSuccess_894);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_895", put_index_895);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_896", put_size_896);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_897", put_isLeaf_897);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_898", put_nextFree_898);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_899", put_Key_0_899);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_900", put_KeyCompares_0_900);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_901", put_KeyCollapse_0_901);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_902", put_Data_0_902);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_903", put_Key_1_903);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_904", put_KeyCompares_1_904);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_905", put_KeyCollapse_1_905);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_906", put_Data_1_906);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_907", put_Key_2_907);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_908", put_KeyCompares_2_908);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_909", put_KeyCollapse_2_909);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_910", put_Data_2_910);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_911", put_Key_3_911);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_912", put_KeyCompares_3_912);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_913", put_KeyCollapse_3_913);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_914", put_Data_3_914);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_915", put_Found_915);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_916", put_Key_916);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_917", put_FoundKey_917);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_918", put_Data_918);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_919", put_BtreeIndex_919);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_920", put_StuckIndex_920);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_921", put_MergeSuccess_921);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_922", put_index_922);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_923", put_size_923);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_924", put_isLeaf_924);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_925", put_nextFree_925);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_926", put_Key_0_926);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_927", put_KeyCompares_0_927);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_928", put_KeyCollapse_0_928);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_929", put_Data_0_929);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_930", put_Key_1_930);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_931", put_KeyCompares_1_931);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_932", put_KeyCollapse_1_932);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_933", put_Data_1_933);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_934", put_Key_2_934);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_935", put_KeyCompares_2_935);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_936", put_KeyCollapse_2_936);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_937", put_Data_2_937);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_938", put_Key_3_938);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_939", put_KeyCompares_3_939);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_940", put_KeyCollapse_3_940);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_941", put_Data_3_941);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_942", put_Found_942);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_943", put_Key_943);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_944", put_FoundKey_944);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_945", put_Data_945);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_946", put_BtreeIndex_946);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_947", put_StuckIndex_947);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_948", put_MergeSuccess_948);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_949", put_childKey_949);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_leftChild_950", put_leftChild_950);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_rightChild_951", put_rightChild_951);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_952", put_childData_952);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_953", put_indexLeft_953);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_954", put_indexRight_954);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_955", put_midKey_955);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_956", put_success_956);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_957", put_test_957);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_958", put_next_958);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_959", put_root_959);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_960", put_isFree_960);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_961", put_next_961);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_962", put_root_962);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_963", put_isFree_963);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_964", put_index_964);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_965", put_size_965);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_966", put_isLeaf_966);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_967", put_nextFree_967);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_968", put_Key_0_968);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_969", put_KeyCompares_0_969);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_970", put_KeyCollapse_0_970);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_971", put_Data_0_971);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_972", put_Key_1_972);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_973", put_KeyCompares_1_973);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_974", put_KeyCollapse_1_974);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_975", put_Data_1_975);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_976", put_Key_2_976);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_977", put_KeyCompares_2_977);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_978", put_KeyCollapse_2_978);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_979", put_Data_2_979);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_980", put_Key_3_980);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_981", put_KeyCompares_3_981);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_982", put_KeyCollapse_3_982);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_983", put_Data_3_983);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_984", put_Found_984);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_985", put_Key_985);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_986", put_FoundKey_986);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_987", put_Data_987);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_988", put_BtreeIndex_988);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_989", put_StuckIndex_989);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_990", put_MergeSuccess_990);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_991", put_index_991);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_992", put_size_992);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_993", put_isLeaf_993);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_994", put_nextFree_994);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_995", put_Key_0_995);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_996", put_KeyCompares_0_996);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_997", put_KeyCollapse_0_997);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_998", put_Data_0_998);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_999", put_Key_1_999);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1000", put_KeyCompares_1_1000);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1001", put_KeyCollapse_1_1001);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1002", put_Data_1_1002);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1003", put_Key_2_1003);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1004", put_KeyCompares_2_1004);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1005", put_KeyCollapse_2_1005);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1006", put_Data_2_1006);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1007", put_Key_3_1007);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1008", put_KeyCompares_3_1008);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1009", put_KeyCollapse_3_1009);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1010", put_Data_3_1010);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1011", put_Found_1011);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1012", put_Key_1012);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1013", put_FoundKey_1013);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1014", put_Data_1014);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1015", put_BtreeIndex_1015);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1016", put_StuckIndex_1016);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1017", put_MergeSuccess_1017);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1018", put_childKey_1018);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1019", put_size_1019);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1020", put_childData_1020);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1021", put_indexLeft_1021);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1022", put_indexRight_1022);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1023", put_midKey_1023);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1024", put_success_1024);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1025", put_test_1025);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1026", put_next_1026);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1027", put_root_1027);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1028", put_isFree_1028);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1029", put_index_1029);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1030", put_size_1030);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1031", put_isLeaf_1031);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1032", put_nextFree_1032);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1033", put_Key_0_1033);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1034", put_KeyCompares_0_1034);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1035", put_KeyCollapse_0_1035);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1036", put_Data_0_1036);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1037", put_Key_1_1037);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1038", put_KeyCompares_1_1038);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1039", put_KeyCollapse_1_1039);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1040", put_Data_1_1040);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1041", put_Key_2_1041);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1042", put_KeyCompares_2_1042);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1043", put_KeyCollapse_2_1043);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1044", put_Data_2_1044);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1045", put_Key_3_1045);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1046", put_KeyCompares_3_1046);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1047", put_KeyCollapse_3_1047);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1048", put_Data_3_1048);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1049", put_Found_1049);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1050", put_Key_1050);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1051", put_FoundKey_1051);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1052", put_Data_1052);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1053", put_BtreeIndex_1053);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1054", put_StuckIndex_1054);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1055", put_MergeSuccess_1055);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1056", put_index_1056);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1057", put_size_1057);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1058", put_isLeaf_1058);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1059", put_nextFree_1059);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1060", put_Key_0_1060);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1061", put_KeyCompares_0_1061);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1062", put_KeyCollapse_0_1062);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1063", put_Data_0_1063);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1064", put_Key_1_1064);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1065", put_KeyCompares_1_1065);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1066", put_KeyCollapse_1_1066);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1067", put_Data_1_1067);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1068", put_Key_2_1068);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1069", put_KeyCompares_2_1069);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1070", put_KeyCollapse_2_1070);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1071", put_Data_2_1071);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1072", put_Key_3_1072);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1073", put_KeyCompares_3_1073);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1074", put_KeyCollapse_3_1074);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1075", put_Data_3_1075);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1076", put_Found_1076);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1077", put_Key_1077);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1078", put_FoundKey_1078);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1079", put_Data_1079);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1080", put_BtreeIndex_1080);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1081", put_StuckIndex_1081);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1082", put_MergeSuccess_1082);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1083", put_childKey_1083);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1084", put_size_1084);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1085", put_childData_1085);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1086", put_indexLeft_1086);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1087", put_indexRight_1087);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1088", put_midKey_1088);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1089", put_success_1089);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1090", put_test_1090);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1091", put_next_1091);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1092", put_root_1092);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1093", put_isFree_1093);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1094", put_index_1094);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1095", put_size_1095);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1096", put_isLeaf_1096);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1097", put_nextFree_1097);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1098", put_Key_0_1098);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1099", put_KeyCompares_0_1099);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1100", put_KeyCollapse_0_1100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1101", put_Data_0_1101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1102", put_Key_1_1102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1103", put_KeyCompares_1_1103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1104", put_KeyCollapse_1_1104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1105", put_Data_1_1105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1106", put_Key_2_1106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1107", put_KeyCompares_2_1107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1108", put_KeyCollapse_2_1108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1109", put_Data_2_1109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1110", put_Key_3_1110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1111", put_KeyCompares_3_1111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1112", put_KeyCollapse_3_1112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1113", put_Data_3_1113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1114", put_Found_1114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1115", put_Key_1115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1116", put_FoundKey_1116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1117", put_Data_1117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1118", put_BtreeIndex_1118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1119", put_StuckIndex_1119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1120", put_MergeSuccess_1120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1121", put_index_1121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1122", put_size_1122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1123", put_isLeaf_1123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1124", put_nextFree_1124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1125", put_Key_0_1125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1126", put_KeyCompares_0_1126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1127", put_KeyCollapse_0_1127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1128", put_Data_0_1128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1129", put_Key_1_1129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1130", put_KeyCompares_1_1130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1131", put_KeyCollapse_1_1131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1132", put_Data_1_1132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1133", put_Key_2_1133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1134", put_KeyCompares_2_1134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1135", put_KeyCollapse_2_1135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1136", put_Data_2_1136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1137", put_Key_3_1137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1138", put_KeyCompares_3_1138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1139", put_KeyCollapse_3_1139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1140", put_Data_3_1140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1141", put_Found_1141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1142", put_Key_1142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1143", put_FoundKey_1143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1144", put_Data_1144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1145", put_BtreeIndex_1145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1146", put_StuckIndex_1146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1147", put_MergeSuccess_1147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1148", put_childKey_1148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1149", put_childData_1149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1150", put_indexLeft_1150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1151", put_indexRight_1151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1152", put_midKey_1152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1153", put_success_1153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1154", put_test_1154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1155", put_next_1155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1156", put_root_1156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1157", put_isFree_1157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1158", put_index_1158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1159", put_size_1159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1160", put_isLeaf_1160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1161", put_nextFree_1161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1162", put_Key_0_1162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1163", put_KeyCompares_0_1163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1164", put_KeyCollapse_0_1164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1165", put_Data_0_1165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1166", put_Key_1_1166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1167", put_KeyCompares_1_1167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1168", put_KeyCollapse_1_1168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1169", put_Data_1_1169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1170", put_Key_2_1170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1171", put_KeyCompares_2_1171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1172", put_KeyCollapse_2_1172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1173", put_Data_2_1173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1174", put_Key_3_1174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1175", put_KeyCompares_3_1175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1176", put_KeyCollapse_3_1176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1177", put_Data_3_1177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1178", put_Found_1178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1179", put_Key_1179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1180", put_FoundKey_1180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1181", put_Data_1181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1182", put_BtreeIndex_1182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1183", put_StuckIndex_1183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1184", put_MergeSuccess_1184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1185", put_index_1185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1186", put_size_1186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1187", put_isLeaf_1187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1188", put_nextFree_1188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1189", put_Key_0_1189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1190", put_KeyCompares_0_1190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1191", put_KeyCollapse_0_1191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1192", put_Data_0_1192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1193", put_Key_1_1193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1194", put_KeyCompares_1_1194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1195", put_KeyCollapse_1_1195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1196", put_Data_1_1196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1197", put_Key_2_1197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1198", put_KeyCompares_2_1198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1199", put_KeyCollapse_2_1199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1200", put_Data_2_1200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1201", put_Key_3_1201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1202", put_KeyCompares_3_1202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1203", put_KeyCollapse_3_1203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1204", put_Data_3_1204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1205", put_Found_1205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1206", put_Key_1206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1207", put_FoundKey_1207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1208", put_Data_1208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1209", put_BtreeIndex_1209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1210", put_StuckIndex_1210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1211", put_MergeSuccess_1211);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1212", put_childKey_1212);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_leftChild_1213", put_leftChild_1213);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_rightChild_1214", put_rightChild_1214);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1215", put_childData_1215);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1216", put_indexLeft_1216);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1217", put_indexRight_1217);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1218", put_midKey_1218);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1219", put_success_1219);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1220", put_test_1220);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1221", put_next_1221);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1222", put_root_1222);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1223", put_isFree_1223);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1224", put_index_1224);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1225", put_size_1225);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1226", put_isLeaf_1226);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1227", put_nextFree_1227);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1228", put_Key_0_1228);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1229", put_KeyCompares_0_1229);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1230", put_KeyCollapse_0_1230);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1231", put_Data_0_1231);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1232", put_Key_1_1232);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1233", put_KeyCompares_1_1233);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1234", put_KeyCollapse_1_1234);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1235", put_Data_1_1235);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1236", put_Key_2_1236);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1237", put_KeyCompares_2_1237);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1238", put_KeyCollapse_2_1238);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1239", put_Data_2_1239);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1240", put_Key_3_1240);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1241", put_KeyCompares_3_1241);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1242", put_KeyCollapse_3_1242);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1243", put_Data_3_1243);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1244", put_Found_1244);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1245", put_Key_1245);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1246", put_FoundKey_1246);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1247", put_Data_1247);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1248", put_BtreeIndex_1248);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1249", put_StuckIndex_1249);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1250", put_MergeSuccess_1250);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1251", put_index_1251);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1252", put_size_1252);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1253", put_isLeaf_1253);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1254", put_nextFree_1254);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1255", put_Key_0_1255);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1256", put_KeyCompares_0_1256);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1257", put_KeyCollapse_0_1257);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1258", put_Data_0_1258);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1259", put_Key_1_1259);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1260", put_KeyCompares_1_1260);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1261", put_KeyCollapse_1_1261);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1262", put_Data_1_1262);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1263", put_Key_2_1263);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1264", put_KeyCompares_2_1264);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1265", put_KeyCollapse_2_1265);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1266", put_Data_2_1266);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1267", put_Key_3_1267);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1268", put_KeyCompares_3_1268);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1269", put_KeyCollapse_3_1269);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1270", put_Data_3_1270);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1271", put_Found_1271);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1272", put_Key_1272);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1273", put_FoundKey_1273);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1274", put_Data_1274);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1275", put_BtreeIndex_1275);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1276", put_StuckIndex_1276);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1277", put_MergeSuccess_1277);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1278", put_childKey_1278);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1279", put_childData_1279);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1280", put_indexLeft_1280);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1281", put_indexRight_1281);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1282", put_midKey_1282);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1283", put_success_1283);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1284", put_test_1284);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1285", put_next_1285);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1286", put_root_1286);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1287", put_isFree_1287);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1288", put_index_1288);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1289", put_size_1289);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1290", put_isLeaf_1290);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1291", put_nextFree_1291);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1292", put_Key_0_1292);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1293", put_KeyCompares_0_1293);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1294", put_KeyCollapse_0_1294);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1295", put_Data_0_1295);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1296", put_Key_1_1296);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1297", put_KeyCompares_1_1297);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1298", put_KeyCollapse_1_1298);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1299", put_Data_1_1299);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1300", put_Key_2_1300);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1301", put_KeyCompares_2_1301);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1302", put_KeyCollapse_2_1302);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1303", put_Data_2_1303);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1304", put_Key_3_1304);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1305", put_KeyCompares_3_1305);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1306", put_KeyCollapse_3_1306);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1307", put_Data_3_1307);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1308", put_Found_1308);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1309", put_Key_1309);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1310", put_FoundKey_1310);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1311", put_Data_1311);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1312", put_BtreeIndex_1312);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1313", put_StuckIndex_1313);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1314", put_MergeSuccess_1314);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1315", put_index_1315);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1316", put_size_1316);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1317", put_isLeaf_1317);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1318", put_nextFree_1318);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1319", put_Key_0_1319);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1320", put_KeyCompares_0_1320);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1321", put_KeyCollapse_0_1321);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1322", put_Data_0_1322);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1323", put_Key_1_1323);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1324", put_KeyCompares_1_1324);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1325", put_KeyCollapse_1_1325);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1326", put_Data_1_1326);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1327", put_Key_2_1327);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1328", put_KeyCompares_2_1328);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1329", put_KeyCollapse_2_1329);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1330", put_Data_2_1330);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1331", put_Key_3_1331);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1332", put_KeyCompares_3_1332);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1333", put_KeyCollapse_3_1333);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1334", put_Data_3_1334);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1335", put_Found_1335);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1336", put_Key_1336);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1337", put_FoundKey_1337);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1338", put_Data_1338);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1339", put_BtreeIndex_1339);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1340", put_StuckIndex_1340);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1341", put_MergeSuccess_1341);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1342", put_childKey_1342);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_leftChild_1343", put_leftChild_1343);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_rightChild_1344", put_rightChild_1344);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1345", put_childData_1345);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1346", put_indexLeft_1346);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1347", put_indexRight_1347);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1348", put_midKey_1348);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1349", put_success_1349);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1350", put_test_1350);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1351", put_next_1351);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1352", put_root_1352);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1353", put_isFree_1353);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1354", put_index_1354);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1355", put_size_1355);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1356", put_isLeaf_1356);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1357", put_nextFree_1357);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1358", put_Key_0_1358);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1359", put_KeyCompares_0_1359);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1360", put_KeyCollapse_0_1360);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1361", put_Data_0_1361);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1362", put_Key_1_1362);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1363", put_KeyCompares_1_1363);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1364", put_KeyCollapse_1_1364);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1365", put_Data_1_1365);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1366", put_Key_2_1366);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1367", put_KeyCompares_2_1367);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1368", put_KeyCollapse_2_1368);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1369", put_Data_2_1369);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1370", put_Key_3_1370);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1371", put_KeyCompares_3_1371);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1372", put_KeyCollapse_3_1372);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1373", put_Data_3_1373);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1374", put_Found_1374);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1375", put_Key_1375);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1376", put_FoundKey_1376);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1377", put_Data_1377);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1378", put_BtreeIndex_1378);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1379", put_StuckIndex_1379);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1380", put_MergeSuccess_1380);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1381", put_index_1381);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1382", put_size_1382);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1383", put_isLeaf_1383);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1384", put_nextFree_1384);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1385", put_Key_0_1385);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1386", put_KeyCompares_0_1386);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1387", put_KeyCollapse_0_1387);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1388", put_Data_0_1388);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1389", put_Key_1_1389);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1390", put_KeyCompares_1_1390);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1391", put_KeyCollapse_1_1391);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1392", put_Data_1_1392);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1393", put_Key_2_1393);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1394", put_KeyCompares_2_1394);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1395", put_KeyCollapse_2_1395);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1396", put_Data_2_1396);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1397", put_Key_3_1397);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1398", put_KeyCompares_3_1398);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1399", put_KeyCollapse_3_1399);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1400", put_Data_3_1400);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1401", put_Found_1401);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1402", put_Key_1402);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1403", put_FoundKey_1403);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1404", put_Data_1404);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1405", put_BtreeIndex_1405);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1406", put_StuckIndex_1406);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1407", put_MergeSuccess_1407);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1408", put_childKey_1408);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1409", put_childData_1409);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1410", put_indexLeft_1410);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1411", put_indexRight_1411);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1412", put_midKey_1412);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1413", put_success_1413);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1414", put_test_1414);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1415", put_next_1415);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1416", put_root_1416);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1417", put_isFree_1417);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1418", put_index_1418);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1419", put_size_1419);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1420", put_isLeaf_1420);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1421", put_nextFree_1421);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1422", put_Key_0_1422);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1423", put_KeyCompares_0_1423);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1424", put_KeyCollapse_0_1424);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1425", put_Data_0_1425);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1426", put_Key_1_1426);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1427", put_KeyCompares_1_1427);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1428", put_KeyCollapse_1_1428);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1429", put_Data_1_1429);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1430", put_Key_2_1430);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1431", put_KeyCompares_2_1431);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1432", put_KeyCollapse_2_1432);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1433", put_Data_2_1433);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1434", put_Key_3_1434);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1435", put_KeyCompares_3_1435);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1436", put_KeyCollapse_3_1436);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1437", put_Data_3_1437);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1438", put_Found_1438);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1439", put_Key_1439);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1440", put_FoundKey_1440);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1441", put_Data_1441);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1442", put_BtreeIndex_1442);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1443", put_StuckIndex_1443);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1444", put_MergeSuccess_1444);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_1445", put_index_1445);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_1446", put_size_1446);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_1447", put_isLeaf_1447);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_1448", put_nextFree_1448);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_1449", put_Key_0_1449);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_1450", put_KeyCompares_0_1450);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_1451", put_KeyCollapse_0_1451);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_1452", put_Data_0_1452);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_1453", put_Key_1_1453);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_1454", put_KeyCompares_1_1454);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_1455", put_KeyCollapse_1_1455);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_1456", put_Data_1_1456);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_1457", put_Key_2_1457);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_1458", put_KeyCompares_2_1458);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_1459", put_KeyCollapse_2_1459);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_1460", put_Data_2_1460);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_1461", put_Key_3_1461);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_1462", put_KeyCompares_3_1462);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_1463", put_KeyCollapse_3_1463);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_1464", put_Data_3_1464);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_1465", put_Found_1465);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1466", put_Key_1466);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_1467", put_FoundKey_1467);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1468", put_Data_1468);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_1469", put_BtreeIndex_1469);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_1470", put_StuckIndex_1470);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_1471", put_MergeSuccess_1471);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_1472", put_childKey_1472);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_leftChild_1473", put_leftChild_1473);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_rightChild_1474", put_rightChild_1474);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_1475", put_childData_1475);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_1476", put_indexLeft_1476);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_1477", put_indexRight_1477);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_1478", put_midKey_1478);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_success_1479", put_success_1479);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_test_1480", put_test_1480);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_1481", put_next_1481);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_1482", put_root_1482);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_1483", put_isFree_1483);
      $fclose(o);
    end
  endtask
endmodule
