//-----------------------------------------------------------------------------
// Database on a chip synthesis
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree(                                                                      // Test bench for database on a chip
  input                 clock,                                                  // Clock
  input                 reset,                                                  // Reset chip

  input wire [64-1:0] k,
  input wire [64-1:0] d,
  output wire            stop                                            // Program has stopped when this goes high
  );
  integer step;
  integer returnCode;
  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_stop||stuckData_stop||verilogPut_stop;
  always @ (posedge clock) begin
    if (reset) begin
      step <= -2;
    end
    else begin
      step <= step + 1;
    end
  end
  // process_stuckIsLeaf_0000
  // process_stuckIsFree_0001
  // process_freeNext_0002
  // process_stuckSize_0003
  // process_stuckKeys_0004
  // process_stuckData_0005
  // process_verilogPut_0006
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[8*1];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_7_result_0;
  integer stuckIsLeaf_7_requestedAt;
  integer stuckIsLeaf_7_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_7_returnCode;
  integer stuckIsLeaf_8_requestedAt;
  integer stuckIsLeaf_8_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_8_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_7_result_0 <= 0;
      stuckIsLeaf_7_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_7_returnCode <= 0;
      stuckIsLeaf_8_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_8_returnCode <= 0;
      stuckIsLeaf_memory[0] <= 1;
      stuckIsLeaf_memory[1] <= 0;
      stuckIsLeaf_memory[2] <= 0;
      stuckIsLeaf_memory[3] <= 0;
      stuckIsLeaf_memory[4] <= 0;
      stuckIsLeaf_memory[5] <= 0;
      stuckIsLeaf_memory[6] <= 0;
      stuckIsLeaf_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_7_result_0 <= stuckIsLeaf_memory[verilogPut_stuckIsLeaf_7_index_37*1+0];
            stuckIsLeaf_7_finishedAt <= step;
          end
          else if ((stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step)) begin
            stuckIsLeaf_memory[verilogPut_stuckIsLeaf_8_index_38*1+0] <= verilogPut_stuckIsLeaf_8_value_39;
            stuckIsLeaf_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[8*1];
  integer stuckIsFree_11_requestedAt;
  integer stuckIsFree_11_finishedAt;
  integer stuckIsFree_stuckIsFree_11_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_11_finishedAt <= -1;
      stuckIsFree_stuckIsFree_11_returnCode <= 0;
      stuckIsFree_memory[0] <= 0;
      stuckIsFree_memory[1] <= 1;
      stuckIsFree_memory[2] <= 1;
      stuckIsFree_memory[3] <= 1;
      stuckIsFree_memory[4] <= 1;
      stuckIsFree_memory[5] <= 1;
      stuckIsFree_memory[6] <= 1;
      stuckIsFree_memory[7] <= 1;
    end
    else begin                                   // Run the process in full parallel
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step)) begin
            stuckIsFree_memory[verilogPut_stuckIsFree_11_index_195*1+0] <= verilogPut_stuckIsFree_11_value_196;
            stuckIsFree_11_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [4-1:0] freeNext_memory[8*1];
  reg [4-1:0] freeNext_freeNext_9_result_0;
  integer freeNext_9_requestedAt;
  integer freeNext_9_finishedAt;
  integer freeNext_freeNext_9_returnCode;
  integer freeNext_10_requestedAt;
  integer freeNext_10_finishedAt;
  integer freeNext_freeNext_10_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_9_result_0 <= 0;
      freeNext_9_finishedAt <= -1;
      freeNext_freeNext_9_returnCode <= 0;
      freeNext_10_finishedAt <= -1;
      freeNext_freeNext_10_returnCode <= 0;
      freeNext_memory[0] <= 1;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 7;
      freeNext_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(freeNext_pc)
        0: begin
          if ((freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step)) begin
            freeNext_freeNext_9_result_0 <= freeNext_memory[verilogPut_freeNext_9_index_192*1+0];
            freeNext_9_finishedAt <= step;
          end
          else if ((freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step)) begin
            freeNext_memory[verilogPut_freeNext_10_index_193*1+0] <= verilogPut_freeNext_10_value_194;
            freeNext_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[8*1];
  reg [3-1:0] stuckSize_stuckSize_5_result_0;
  integer stuckSize_5_requestedAt;
  integer stuckSize_5_finishedAt;
  integer stuckSize_stuckSize_5_returnCode;
  integer stuckSize_6_requestedAt;
  integer stuckSize_6_finishedAt;
  integer stuckSize_stuckSize_6_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_5_result_0 <= 0;
      stuckSize_5_finishedAt <= -1;
      stuckSize_stuckSize_5_returnCode <= 0;
      stuckSize_6_finishedAt <= -1;
      stuckSize_stuckSize_6_returnCode <= 0;
      stuckSize_memory[0] <= 0;
      stuckSize_memory[1] <= 0;
      stuckSize_memory[2] <= 0;
      stuckSize_memory[3] <= 0;
      stuckSize_memory[4] <= 0;
      stuckSize_memory[5] <= 0;
      stuckSize_memory[6] <= 0;
      stuckSize_memory[7] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step)) begin
            stuckSize_stuckSize_5_result_0 <= stuckSize_memory[verilogPut_stuckSize_5_index_34*1+0];
            stuckSize_5_finishedAt <= step;
          end
          else if ((stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step)) begin
            stuckSize_memory[verilogPut_stuckSize_6_index_35*1+0] <= verilogPut_stuckSize_6_value_36;
            stuckSize_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys  process_stuckKeys_0004
  (* ram_style = "block" *)
  reg [64-1:0] stuckKeys_memory[8*4];
  reg [64-1:0] stuckKeys_stuckKeys_1_result_0;
  reg [64-1:0] stuckKeys_stuckKeys_1_result_1;
  reg [64-1:0] stuckKeys_stuckKeys_1_result_2;
  reg [64-1:0] stuckKeys_stuckKeys_1_result_3;
  integer stuckKeys_1_requestedAt;
  integer stuckKeys_1_finishedAt;
  integer stuckKeys_stuckKeys_1_returnCode;
  integer stuckKeys_2_requestedAt;
  integer stuckKeys_2_finishedAt;
  integer stuckKeys_stuckKeys_2_returnCode;
  integer stuckKeys_pc;
  integer stuckKeys_stop;
  integer stuckKeys_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_pc <= 0;
      stuckKeys_stop <= 0;
      stuckKeys_returnCode <= 0;
      stuckKeys_stuckKeys_1_result_0 <= 0;
      stuckKeys_stuckKeys_1_result_1 <= 0;
      stuckKeys_stuckKeys_1_result_2 <= 0;
      stuckKeys_stuckKeys_1_result_3 <= 0;
      stuckKeys_1_finishedAt <= -1;
      stuckKeys_stuckKeys_1_returnCode <= 0;
      stuckKeys_2_finishedAt <= -1;
      stuckKeys_stuckKeys_2_returnCode <= 0;
      stuckKeys_memory[0] <= 0;
      stuckKeys_memory[1] <= 0;
      stuckKeys_memory[2] <= 0;
      stuckKeys_memory[3] <= 0;
      stuckKeys_memory[4] <= 0;
      stuckKeys_memory[5] <= 0;
      stuckKeys_memory[6] <= 0;
      stuckKeys_memory[7] <= 0;
      stuckKeys_memory[8] <= 0;
      stuckKeys_memory[9] <= 0;
      stuckKeys_memory[10] <= 0;
      stuckKeys_memory[11] <= 0;
      stuckKeys_memory[12] <= 0;
      stuckKeys_memory[13] <= 0;
      stuckKeys_memory[14] <= 0;
      stuckKeys_memory[15] <= 0;
      stuckKeys_memory[16] <= 0;
      stuckKeys_memory[17] <= 0;
      stuckKeys_memory[18] <= 0;
      stuckKeys_memory[19] <= 0;
      stuckKeys_memory[20] <= 0;
      stuckKeys_memory[21] <= 0;
      stuckKeys_memory[22] <= 0;
      stuckKeys_memory[23] <= 0;
      stuckKeys_memory[24] <= 0;
      stuckKeys_memory[25] <= 0;
      stuckKeys_memory[26] <= 0;
      stuckKeys_memory[27] <= 0;
      stuckKeys_memory[28] <= 0;
      stuckKeys_memory[29] <= 0;
      stuckKeys_memory[30] <= 0;
      stuckKeys_memory[31] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckKeys_pc)
        0: begin
          if ((stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step)) begin
            stuckKeys_stuckKeys_1_result_0 <= stuckKeys_memory[verilogPut_stuckKeys_1_index_22*4+0];
            stuckKeys_stuckKeys_1_result_1 <= stuckKeys_memory[verilogPut_stuckKeys_1_index_22*4+1];
            stuckKeys_stuckKeys_1_result_2 <= stuckKeys_memory[verilogPut_stuckKeys_1_index_22*4+2];
            stuckKeys_stuckKeys_1_result_3 <= stuckKeys_memory[verilogPut_stuckKeys_1_index_22*4+3];
            stuckKeys_1_finishedAt <= step;
          end
          else if ((stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step)) begin
            stuckKeys_memory[verilogPut_stuckKeys_2_index_23*4+0] <= verilogPut_stuckKeys_2_value_24;
            stuckKeys_memory[verilogPut_stuckKeys_2_index_23*4+1] <= verilogPut_stuckKeys_2_value_25;
            stuckKeys_memory[verilogPut_stuckKeys_2_index_23*4+2] <= verilogPut_stuckKeys_2_value_26;
            stuckKeys_memory[verilogPut_stuckKeys_2_index_23*4+3] <= verilogPut_stuckKeys_2_value_27;
            stuckKeys_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_stop <= 1;
      endcase
    end
  end
  // Process: stuckData  process_stuckData_0005
  (* ram_style = "block" *)
  reg [64-1:0] stuckData_memory[8*4];
  reg [64-1:0] stuckData_stuckData_3_result_0;
  reg [64-1:0] stuckData_stuckData_3_result_1;
  reg [64-1:0] stuckData_stuckData_3_result_2;
  reg [64-1:0] stuckData_stuckData_3_result_3;
  integer stuckData_3_requestedAt;
  integer stuckData_3_finishedAt;
  integer stuckData_stuckData_3_returnCode;
  integer stuckData_4_requestedAt;
  integer stuckData_4_finishedAt;
  integer stuckData_stuckData_4_returnCode;
  integer stuckData_pc;
  integer stuckData_stop;
  integer stuckData_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_pc <= 0;
      stuckData_stop <= 0;
      stuckData_returnCode <= 0;
      stuckData_stuckData_3_result_0 <= 0;
      stuckData_stuckData_3_result_1 <= 0;
      stuckData_stuckData_3_result_2 <= 0;
      stuckData_stuckData_3_result_3 <= 0;
      stuckData_3_finishedAt <= -1;
      stuckData_stuckData_3_returnCode <= 0;
      stuckData_4_finishedAt <= -1;
      stuckData_stuckData_4_returnCode <= 0;
      stuckData_memory[0] <= 0;
      stuckData_memory[1] <= 0;
      stuckData_memory[2] <= 0;
      stuckData_memory[3] <= 0;
      stuckData_memory[4] <= 0;
      stuckData_memory[5] <= 0;
      stuckData_memory[6] <= 0;
      stuckData_memory[7] <= 0;
      stuckData_memory[8] <= 0;
      stuckData_memory[9] <= 0;
      stuckData_memory[10] <= 0;
      stuckData_memory[11] <= 0;
      stuckData_memory[12] <= 0;
      stuckData_memory[13] <= 0;
      stuckData_memory[14] <= 0;
      stuckData_memory[15] <= 0;
      stuckData_memory[16] <= 0;
      stuckData_memory[17] <= 0;
      stuckData_memory[18] <= 0;
      stuckData_memory[19] <= 0;
      stuckData_memory[20] <= 0;
      stuckData_memory[21] <= 0;
      stuckData_memory[22] <= 0;
      stuckData_memory[23] <= 0;
      stuckData_memory[24] <= 0;
      stuckData_memory[25] <= 0;
      stuckData_memory[26] <= 0;
      stuckData_memory[27] <= 0;
      stuckData_memory[28] <= 0;
      stuckData_memory[29] <= 0;
      stuckData_memory[30] <= 0;
      stuckData_memory[31] <= 0;
    end
    else begin                                   // Run the process in full parallel
      case(stuckData_pc)
        0: begin
          if ((stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step)) begin
            stuckData_stuckData_3_result_0 <= stuckData_memory[verilogPut_stuckData_3_index_28*4+0];
            stuckData_stuckData_3_result_1 <= stuckData_memory[verilogPut_stuckData_3_index_28*4+1];
            stuckData_stuckData_3_result_2 <= stuckData_memory[verilogPut_stuckData_3_index_28*4+2];
            stuckData_stuckData_3_result_3 <= stuckData_memory[verilogPut_stuckData_3_index_28*4+3];
            stuckData_3_finishedAt <= step;
          end
          else if ((stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step)) begin
            stuckData_memory[verilogPut_stuckData_4_index_29*4+0] <= verilogPut_stuckData_4_value_30;
            stuckData_memory[verilogPut_stuckData_4_index_29*4+1] <= verilogPut_stuckData_4_value_31;
            stuckData_memory[verilogPut_stuckData_4_index_29*4+2] <= verilogPut_stuckData_4_value_32;
            stuckData_memory[verilogPut_stuckData_4_index_29*4+3] <= verilogPut_stuckData_4_value_33;
            stuckData_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_stop <= 1;
      endcase
    end
  end
  // Process: verilogPut  process_verilogPut_0006
  reg [64-1:0] verilogPut_k_0;
  reg [64-1:0] verilogPut_d_1;
  reg [4-1:0] verilogPut_index_2;
  reg [3-1:0] verilogPut_size_3;
  reg [1-1:0] verilogPut_isLeaf_4;
  reg [4-1:0] verilogPut_nextFree_5;
  reg [64-1:0] verilogPut_Key_0_6;
  reg [1-1:0] verilogPut_KeyCompares_0_7;
  reg [3-1:0] verilogPut_KeyCollapse_0_8;
  reg [64-1:0] verilogPut_Data_0_9;
  reg [64-1:0] verilogPut_Key_1_10;
  reg [1-1:0] verilogPut_KeyCompares_1_11;
  reg [3-1:0] verilogPut_KeyCollapse_1_12;
  reg [64-1:0] verilogPut_Data_1_13;
  reg [64-1:0] verilogPut_Key_2_14;
  reg [1-1:0] verilogPut_KeyCompares_2_15;
  reg [3-1:0] verilogPut_KeyCollapse_2_16;
  reg [64-1:0] verilogPut_Data_2_17;
  reg [64-1:0] verilogPut_Key_3_18;
  reg [1-1:0] verilogPut_KeyCompares_3_19;
  reg [3-1:0] verilogPut_KeyCollapse_3_20;
  reg [64-1:0] verilogPut_Data_3_21;
  reg [3-1:0] verilogPut_stuckKeys_1_index_22;
  reg [3-1:0] verilogPut_stuckKeys_2_index_23;
  reg [64-1:0] verilogPut_stuckKeys_2_value_24;
  reg [64-1:0] verilogPut_stuckKeys_2_value_25;
  reg [64-1:0] verilogPut_stuckKeys_2_value_26;
  reg [64-1:0] verilogPut_stuckKeys_2_value_27;
  reg [3-1:0] verilogPut_stuckData_3_index_28;
  reg [3-1:0] verilogPut_stuckData_4_index_29;
  reg [64-1:0] verilogPut_stuckData_4_value_30;
  reg [64-1:0] verilogPut_stuckData_4_value_31;
  reg [64-1:0] verilogPut_stuckData_4_value_32;
  reg [64-1:0] verilogPut_stuckData_4_value_33;
  reg [3-1:0] verilogPut_stuckSize_5_index_34;
  reg [3-1:0] verilogPut_stuckSize_6_index_35;
  reg [3-1:0] verilogPut_stuckSize_6_value_36;
  reg [3-1:0] verilogPut_stuckIsLeaf_7_index_37;
  reg [3-1:0] verilogPut_stuckIsLeaf_8_index_38;
  reg [1-1:0] verilogPut_stuckIsLeaf_8_value_39;
  reg [1-1:0] verilogPut_Found_40;
  reg [64-1:0] verilogPut_Key_41;
  reg [64-1:0] verilogPut_FoundKey_42;
  reg [64-1:0] verilogPut_Data_43;
  reg [4-1:0] verilogPut_BtreeIndex_44;
  reg [3-1:0] verilogPut_StuckIndex_45;
  reg [1-1:0] verilogPut_MergeSuccess_46;
  reg [4-1:0] verilogPut_index_47;
  reg [3-1:0] verilogPut_size_48;
  reg [1-1:0] verilogPut_isLeaf_49;
  reg [4-1:0] verilogPut_nextFree_50;
  reg [64-1:0] verilogPut_Key_0_51;
  reg [1-1:0] verilogPut_KeyCompares_0_52;
  reg [3-1:0] verilogPut_KeyCollapse_0_53;
  reg [64-1:0] verilogPut_Data_0_54;
  reg [64-1:0] verilogPut_Key_1_55;
  reg [1-1:0] verilogPut_KeyCompares_1_56;
  reg [3-1:0] verilogPut_KeyCollapse_1_57;
  reg [64-1:0] verilogPut_Data_1_58;
  reg [64-1:0] verilogPut_Key_2_59;
  reg [1-1:0] verilogPut_KeyCompares_2_60;
  reg [3-1:0] verilogPut_KeyCollapse_2_61;
  reg [64-1:0] verilogPut_Data_2_62;
  reg [64-1:0] verilogPut_Key_3_63;
  reg [1-1:0] verilogPut_KeyCompares_3_64;
  reg [3-1:0] verilogPut_KeyCollapse_3_65;
  reg [64-1:0] verilogPut_Data_3_66;
  reg [1-1:0] verilogPut_Found_67;
  reg [64-1:0] verilogPut_Key_68;
  reg [64-1:0] verilogPut_FoundKey_69;
  reg [64-1:0] verilogPut_Data_70;
  reg [4-1:0] verilogPut_BtreeIndex_71;
  reg [3-1:0] verilogPut_StuckIndex_72;
  reg [1-1:0] verilogPut_MergeSuccess_73;
  reg [4-1:0] verilogPut_index_74;
  reg [3-1:0] verilogPut_size_75;
  reg [1-1:0] verilogPut_isLeaf_76;
  reg [4-1:0] verilogPut_nextFree_77;
  reg [64-1:0] verilogPut_Key_0_78;
  reg [1-1:0] verilogPut_KeyCompares_0_79;
  reg [3-1:0] verilogPut_KeyCollapse_0_80;
  reg [64-1:0] verilogPut_Data_0_81;
  reg [64-1:0] verilogPut_Key_1_82;
  reg [1-1:0] verilogPut_KeyCompares_1_83;
  reg [3-1:0] verilogPut_KeyCollapse_1_84;
  reg [64-1:0] verilogPut_Data_1_85;
  reg [64-1:0] verilogPut_Key_2_86;
  reg [1-1:0] verilogPut_KeyCompares_2_87;
  reg [3-1:0] verilogPut_KeyCollapse_2_88;
  reg [64-1:0] verilogPut_Data_2_89;
  reg [64-1:0] verilogPut_Key_3_90;
  reg [1-1:0] verilogPut_KeyCompares_3_91;
  reg [3-1:0] verilogPut_KeyCollapse_3_92;
  reg [64-1:0] verilogPut_Data_3_93;
  reg [1-1:0] verilogPut_Found_94;
  reg [64-1:0] verilogPut_Key_95;
  reg [64-1:0] verilogPut_FoundKey_96;
  reg [64-1:0] verilogPut_Data_97;
  reg [4-1:0] verilogPut_BtreeIndex_98;
  reg [3-1:0] verilogPut_StuckIndex_99;
  reg [1-1:0] verilogPut_MergeSuccess_100;
  reg [4-1:0] verilogPut_child_101;
  reg [4-1:0] verilogPut_parent_102;
  reg [3-1:0] verilogPut_childInparent_103;
  reg [1-1:0] verilogPut_found_104;
  reg [1-1:0] verilogPut_full_105;
  reg [3-1:0] verilogPut_i_106;
  reg [1-1:0] verilogPut_notFull_107;
  reg [4-1:0] verilogPut_index_108;
  reg [3-1:0] verilogPut_size_109;
  reg [1-1:0] verilogPut_isLeaf_110;
  reg [4-1:0] verilogPut_nextFree_111;
  reg [64-1:0] verilogPut_Key_0_112;
  reg [1-1:0] verilogPut_KeyCompares_0_113;
  reg [3-1:0] verilogPut_KeyCollapse_0_114;
  reg [64-1:0] verilogPut_Data_0_115;
  reg [64-1:0] verilogPut_Key_1_116;
  reg [1-1:0] verilogPut_KeyCompares_1_117;
  reg [3-1:0] verilogPut_KeyCollapse_1_118;
  reg [64-1:0] verilogPut_Data_1_119;
  reg [64-1:0] verilogPut_Key_2_120;
  reg [1-1:0] verilogPut_KeyCompares_2_121;
  reg [3-1:0] verilogPut_KeyCollapse_2_122;
  reg [64-1:0] verilogPut_Data_2_123;
  reg [64-1:0] verilogPut_Key_3_124;
  reg [1-1:0] verilogPut_KeyCompares_3_125;
  reg [3-1:0] verilogPut_KeyCollapse_3_126;
  reg [64-1:0] verilogPut_Data_3_127;
  reg [1-1:0] verilogPut_Found_128;
  reg [64-1:0] verilogPut_Key_129;
  reg [64-1:0] verilogPut_FoundKey_130;
  reg [64-1:0] verilogPut_Data_131;
  reg [4-1:0] verilogPut_BtreeIndex_132;
  reg [3-1:0] verilogPut_StuckIndex_133;
  reg [1-1:0] verilogPut_MergeSuccess_134;
  reg [4-1:0] verilogPut_index_135;
  reg [3-1:0] verilogPut_size_136;
  reg [1-1:0] verilogPut_isLeaf_137;
  reg [4-1:0] verilogPut_nextFree_138;
  reg [64-1:0] verilogPut_Key_0_139;
  reg [1-1:0] verilogPut_KeyCompares_0_140;
  reg [3-1:0] verilogPut_KeyCollapse_0_141;
  reg [64-1:0] verilogPut_Data_0_142;
  reg [64-1:0] verilogPut_Key_1_143;
  reg [1-1:0] verilogPut_KeyCompares_1_144;
  reg [3-1:0] verilogPut_KeyCollapse_1_145;
  reg [64-1:0] verilogPut_Data_1_146;
  reg [64-1:0] verilogPut_Key_2_147;
  reg [1-1:0] verilogPut_KeyCompares_2_148;
  reg [3-1:0] verilogPut_KeyCollapse_2_149;
  reg [64-1:0] verilogPut_Data_2_150;
  reg [64-1:0] verilogPut_Key_3_151;
  reg [1-1:0] verilogPut_KeyCompares_3_152;
  reg [3-1:0] verilogPut_KeyCollapse_3_153;
  reg [64-1:0] verilogPut_Data_3_154;
  reg [1-1:0] verilogPut_Found_155;
  reg [64-1:0] verilogPut_Key_156;
  reg [64-1:0] verilogPut_FoundKey_157;
  reg [64-1:0] verilogPut_Data_158;
  reg [4-1:0] verilogPut_BtreeIndex_159;
  reg [3-1:0] verilogPut_StuckIndex_160;
  reg [1-1:0] verilogPut_MergeSuccess_161;
  reg [4-1:0] verilogPut_index_162;
  reg [3-1:0] verilogPut_size_163;
  reg [1-1:0] verilogPut_isLeaf_164;
  reg [4-1:0] verilogPut_nextFree_165;
  reg [64-1:0] verilogPut_Key_0_166;
  reg [1-1:0] verilogPut_KeyCompares_0_167;
  reg [3-1:0] verilogPut_KeyCollapse_0_168;
  reg [64-1:0] verilogPut_Data_0_169;
  reg [64-1:0] verilogPut_Key_1_170;
  reg [1-1:0] verilogPut_KeyCompares_1_171;
  reg [3-1:0] verilogPut_KeyCollapse_1_172;
  reg [64-1:0] verilogPut_Data_1_173;
  reg [64-1:0] verilogPut_Key_2_174;
  reg [1-1:0] verilogPut_KeyCompares_2_175;
  reg [3-1:0] verilogPut_KeyCollapse_2_176;
  reg [64-1:0] verilogPut_Data_2_177;
  reg [64-1:0] verilogPut_Key_3_178;
  reg [1-1:0] verilogPut_KeyCompares_3_179;
  reg [3-1:0] verilogPut_KeyCollapse_3_180;
  reg [64-1:0] verilogPut_Data_3_181;
  reg [1-1:0] verilogPut_Found_182;
  reg [64-1:0] verilogPut_Key_183;
  reg [64-1:0] verilogPut_FoundKey_184;
  reg [64-1:0] verilogPut_Data_185;
  reg [4-1:0] verilogPut_BtreeIndex_186;
  reg [3-1:0] verilogPut_StuckIndex_187;
  reg [1-1:0] verilogPut_MergeSuccess_188;
  reg [4-1:0] verilogPut_indexLeft_189;
  reg [4-1:0] verilogPut_indexRight_190;
  reg [64-1:0] verilogPut_midKey_191;
  reg [3-1:0] verilogPut_freeNext_9_index_192;
  reg [3-1:0] verilogPut_freeNext_10_index_193;
  reg [4-1:0] verilogPut_freeNext_10_value_194;
  reg [3-1:0] verilogPut_stuckIsFree_11_index_195;
  reg [1-1:0] verilogPut_stuckIsFree_11_value_196;
  reg [4-1:0] verilogPut_root_197;
  reg [4-1:0] verilogPut_next_198;
  reg [1-1:0] verilogPut_isLeaf_199;
  reg [1-1:0] verilogPut_isFree_200;
  reg [4-1:0] verilogPut_root_201;
  reg [4-1:0] verilogPut_next_202;
  reg [1-1:0] verilogPut_isLeaf_203;
  reg [1-1:0] verilogPut_isFree_204;
  reg [3-1:0] verilogPut_i_205;
  reg [1-1:0] verilogPut_notFull_206;
  reg [4-1:0] verilogPut_index_207;
  reg [3-1:0] verilogPut_size_208;
  reg [1-1:0] verilogPut_isLeaf_209;
  reg [4-1:0] verilogPut_nextFree_210;
  reg [64-1:0] verilogPut_Key_0_211;
  reg [1-1:0] verilogPut_KeyCompares_0_212;
  reg [3-1:0] verilogPut_KeyCollapse_0_213;
  reg [64-1:0] verilogPut_Data_0_214;
  reg [64-1:0] verilogPut_Key_1_215;
  reg [1-1:0] verilogPut_KeyCompares_1_216;
  reg [3-1:0] verilogPut_KeyCollapse_1_217;
  reg [64-1:0] verilogPut_Data_1_218;
  reg [64-1:0] verilogPut_Key_2_219;
  reg [1-1:0] verilogPut_KeyCompares_2_220;
  reg [3-1:0] verilogPut_KeyCollapse_2_221;
  reg [64-1:0] verilogPut_Data_2_222;
  reg [64-1:0] verilogPut_Key_3_223;
  reg [1-1:0] verilogPut_KeyCompares_3_224;
  reg [3-1:0] verilogPut_KeyCollapse_3_225;
  reg [64-1:0] verilogPut_Data_3_226;
  reg [1-1:0] verilogPut_Found_227;
  reg [64-1:0] verilogPut_Key_228;
  reg [64-1:0] verilogPut_FoundKey_229;
  reg [64-1:0] verilogPut_Data_230;
  reg [4-1:0] verilogPut_BtreeIndex_231;
  reg [3-1:0] verilogPut_StuckIndex_232;
  reg [1-1:0] verilogPut_MergeSuccess_233;
  reg [4-1:0] verilogPut_index_234;
  reg [3-1:0] verilogPut_size_235;
  reg [1-1:0] verilogPut_isLeaf_236;
  reg [4-1:0] verilogPut_nextFree_237;
  reg [64-1:0] verilogPut_Key_0_238;
  reg [1-1:0] verilogPut_KeyCompares_0_239;
  reg [3-1:0] verilogPut_KeyCollapse_0_240;
  reg [64-1:0] verilogPut_Data_0_241;
  reg [64-1:0] verilogPut_Key_1_242;
  reg [1-1:0] verilogPut_KeyCompares_1_243;
  reg [3-1:0] verilogPut_KeyCollapse_1_244;
  reg [64-1:0] verilogPut_Data_1_245;
  reg [64-1:0] verilogPut_Key_2_246;
  reg [1-1:0] verilogPut_KeyCompares_2_247;
  reg [3-1:0] verilogPut_KeyCollapse_2_248;
  reg [64-1:0] verilogPut_Data_2_249;
  reg [64-1:0] verilogPut_Key_3_250;
  reg [1-1:0] verilogPut_KeyCompares_3_251;
  reg [3-1:0] verilogPut_KeyCollapse_3_252;
  reg [64-1:0] verilogPut_Data_3_253;
  reg [1-1:0] verilogPut_Found_254;
  reg [64-1:0] verilogPut_Key_255;
  reg [64-1:0] verilogPut_FoundKey_256;
  reg [64-1:0] verilogPut_Data_257;
  reg [4-1:0] verilogPut_BtreeIndex_258;
  reg [3-1:0] verilogPut_StuckIndex_259;
  reg [1-1:0] verilogPut_MergeSuccess_260;
  reg [4-1:0] verilogPut_index_261;
  reg [3-1:0] verilogPut_size_262;
  reg [1-1:0] verilogPut_isLeaf_263;
  reg [4-1:0] verilogPut_nextFree_264;
  reg [64-1:0] verilogPut_Key_0_265;
  reg [1-1:0] verilogPut_KeyCompares_0_266;
  reg [3-1:0] verilogPut_KeyCollapse_0_267;
  reg [64-1:0] verilogPut_Data_0_268;
  reg [64-1:0] verilogPut_Key_1_269;
  reg [1-1:0] verilogPut_KeyCompares_1_270;
  reg [3-1:0] verilogPut_KeyCollapse_1_271;
  reg [64-1:0] verilogPut_Data_1_272;
  reg [64-1:0] verilogPut_Key_2_273;
  reg [1-1:0] verilogPut_KeyCompares_2_274;
  reg [3-1:0] verilogPut_KeyCollapse_2_275;
  reg [64-1:0] verilogPut_Data_2_276;
  reg [64-1:0] verilogPut_Key_3_277;
  reg [1-1:0] verilogPut_KeyCompares_3_278;
  reg [3-1:0] verilogPut_KeyCollapse_3_279;
  reg [64-1:0] verilogPut_Data_3_280;
  reg [1-1:0] verilogPut_Found_281;
  reg [64-1:0] verilogPut_Key_282;
  reg [64-1:0] verilogPut_FoundKey_283;
  reg [64-1:0] verilogPut_Data_284;
  reg [4-1:0] verilogPut_BtreeIndex_285;
  reg [3-1:0] verilogPut_StuckIndex_286;
  reg [1-1:0] verilogPut_MergeSuccess_287;
  reg [4-1:0] verilogPut_indexLeft_288;
  reg [4-1:0] verilogPut_indexRight_289;
  reg [64-1:0] verilogPut_midKey_290;
  reg [4-1:0] verilogPut_root_291;
  reg [4-1:0] verilogPut_next_292;
  reg [1-1:0] verilogPut_isLeaf_293;
  reg [1-1:0] verilogPut_isFree_294;
  reg [4-1:0] verilogPut_root_295;
  reg [4-1:0] verilogPut_next_296;
  reg [1-1:0] verilogPut_isLeaf_297;
  reg [1-1:0] verilogPut_isFree_298;
  reg [4-1:0] verilogPut_index_299;
  reg [3-1:0] verilogPut_size_300;
  reg [1-1:0] verilogPut_isLeaf_301;
  reg [4-1:0] verilogPut_nextFree_302;
  reg [64-1:0] verilogPut_Key_0_303;
  reg [1-1:0] verilogPut_KeyCompares_0_304;
  reg [3-1:0] verilogPut_KeyCollapse_0_305;
  reg [64-1:0] verilogPut_Data_0_306;
  reg [64-1:0] verilogPut_Key_1_307;
  reg [1-1:0] verilogPut_KeyCompares_1_308;
  reg [3-1:0] verilogPut_KeyCollapse_1_309;
  reg [64-1:0] verilogPut_Data_1_310;
  reg [64-1:0] verilogPut_Key_2_311;
  reg [1-1:0] verilogPut_KeyCompares_2_312;
  reg [3-1:0] verilogPut_KeyCollapse_2_313;
  reg [64-1:0] verilogPut_Data_2_314;
  reg [64-1:0] verilogPut_Key_3_315;
  reg [1-1:0] verilogPut_KeyCompares_3_316;
  reg [3-1:0] verilogPut_KeyCollapse_3_317;
  reg [64-1:0] verilogPut_Data_3_318;
  reg [1-1:0] verilogPut_Found_319;
  reg [64-1:0] verilogPut_Key_320;
  reg [64-1:0] verilogPut_FoundKey_321;
  reg [64-1:0] verilogPut_Data_322;
  reg [4-1:0] verilogPut_BtreeIndex_323;
  reg [3-1:0] verilogPut_StuckIndex_324;
  reg [1-1:0] verilogPut_MergeSuccess_325;
  reg [4-1:0] verilogPut_index_326;
  reg [3-1:0] verilogPut_size_327;
  reg [1-1:0] verilogPut_isLeaf_328;
  reg [4-1:0] verilogPut_nextFree_329;
  reg [64-1:0] verilogPut_Key_0_330;
  reg [1-1:0] verilogPut_KeyCompares_0_331;
  reg [3-1:0] verilogPut_KeyCollapse_0_332;
  reg [64-1:0] verilogPut_Data_0_333;
  reg [64-1:0] verilogPut_Key_1_334;
  reg [1-1:0] verilogPut_KeyCompares_1_335;
  reg [3-1:0] verilogPut_KeyCollapse_1_336;
  reg [64-1:0] verilogPut_Data_1_337;
  reg [64-1:0] verilogPut_Key_2_338;
  reg [1-1:0] verilogPut_KeyCompares_2_339;
  reg [3-1:0] verilogPut_KeyCollapse_2_340;
  reg [64-1:0] verilogPut_Data_2_341;
  reg [64-1:0] verilogPut_Key_3_342;
  reg [1-1:0] verilogPut_KeyCompares_3_343;
  reg [3-1:0] verilogPut_KeyCollapse_3_344;
  reg [64-1:0] verilogPut_Data_3_345;
  reg [1-1:0] verilogPut_Found_346;
  reg [64-1:0] verilogPut_Key_347;
  reg [64-1:0] verilogPut_FoundKey_348;
  reg [64-1:0] verilogPut_Data_349;
  reg [4-1:0] verilogPut_BtreeIndex_350;
  reg [3-1:0] verilogPut_StuckIndex_351;
  reg [1-1:0] verilogPut_MergeSuccess_352;
  reg [4-1:0] verilogPut_index_353;
  reg [3-1:0] verilogPut_size_354;
  reg [1-1:0] verilogPut_isLeaf_355;
  reg [4-1:0] verilogPut_nextFree_356;
  reg [64-1:0] verilogPut_Key_0_357;
  reg [1-1:0] verilogPut_KeyCompares_0_358;
  reg [3-1:0] verilogPut_KeyCollapse_0_359;
  reg [64-1:0] verilogPut_Data_0_360;
  reg [64-1:0] verilogPut_Key_1_361;
  reg [1-1:0] verilogPut_KeyCompares_1_362;
  reg [3-1:0] verilogPut_KeyCollapse_1_363;
  reg [64-1:0] verilogPut_Data_1_364;
  reg [64-1:0] verilogPut_Key_2_365;
  reg [1-1:0] verilogPut_KeyCompares_2_366;
  reg [3-1:0] verilogPut_KeyCollapse_2_367;
  reg [64-1:0] verilogPut_Data_2_368;
  reg [64-1:0] verilogPut_Key_3_369;
  reg [1-1:0] verilogPut_KeyCompares_3_370;
  reg [3-1:0] verilogPut_KeyCollapse_3_371;
  reg [64-1:0] verilogPut_Data_3_372;
  reg [1-1:0] verilogPut_Found_373;
  reg [64-1:0] verilogPut_Key_374;
  reg [64-1:0] verilogPut_FoundKey_375;
  reg [64-1:0] verilogPut_Data_376;
  reg [4-1:0] verilogPut_BtreeIndex_377;
  reg [3-1:0] verilogPut_StuckIndex_378;
  reg [1-1:0] verilogPut_MergeSuccess_379;
  reg [4-1:0] verilogPut_index_380;
  reg [3-1:0] verilogPut_size_381;
  reg [1-1:0] verilogPut_isLeaf_382;
  reg [4-1:0] verilogPut_nextFree_383;
  reg [64-1:0] verilogPut_Key_0_384;
  reg [1-1:0] verilogPut_KeyCompares_0_385;
  reg [3-1:0] verilogPut_KeyCollapse_0_386;
  reg [64-1:0] verilogPut_Data_0_387;
  reg [64-1:0] verilogPut_Key_1_388;
  reg [1-1:0] verilogPut_KeyCompares_1_389;
  reg [3-1:0] verilogPut_KeyCollapse_1_390;
  reg [64-1:0] verilogPut_Data_1_391;
  reg [64-1:0] verilogPut_Key_2_392;
  reg [1-1:0] verilogPut_KeyCompares_2_393;
  reg [3-1:0] verilogPut_KeyCollapse_2_394;
  reg [64-1:0] verilogPut_Data_2_395;
  reg [64-1:0] verilogPut_Key_3_396;
  reg [1-1:0] verilogPut_KeyCompares_3_397;
  reg [3-1:0] verilogPut_KeyCollapse_3_398;
  reg [64-1:0] verilogPut_Data_3_399;
  reg [1-1:0] verilogPut_Found_400;
  reg [64-1:0] verilogPut_Key_401;
  reg [64-1:0] verilogPut_FoundKey_402;
  reg [64-1:0] verilogPut_Data_403;
  reg [4-1:0] verilogPut_BtreeIndex_404;
  reg [3-1:0] verilogPut_StuckIndex_405;
  reg [1-1:0] verilogPut_MergeSuccess_406;
  reg [64-1:0] verilogPut_childKey_407;
  reg [4-1:0] verilogPut_childData_408;
  reg [4-1:0] verilogPut_indexLeft_409;
  reg [4-1:0] verilogPut_indexRight_410;
  reg [64-1:0] verilogPut_midKey_411;
  reg [4-1:0] verilogPut_root_412;
  reg [4-1:0] verilogPut_next_413;
  reg [1-1:0] verilogPut_isLeaf_414;
  reg [1-1:0] verilogPut_isFree_415;
  reg [4-1:0] verilogPut_index_416;
  reg [3-1:0] verilogPut_size_417;
  reg [1-1:0] verilogPut_isLeaf_418;
  reg [4-1:0] verilogPut_nextFree_419;
  reg [64-1:0] verilogPut_Key_0_420;
  reg [1-1:0] verilogPut_KeyCompares_0_421;
  reg [3-1:0] verilogPut_KeyCollapse_0_422;
  reg [64-1:0] verilogPut_Data_0_423;
  reg [64-1:0] verilogPut_Key_1_424;
  reg [1-1:0] verilogPut_KeyCompares_1_425;
  reg [3-1:0] verilogPut_KeyCollapse_1_426;
  reg [64-1:0] verilogPut_Data_1_427;
  reg [64-1:0] verilogPut_Key_2_428;
  reg [1-1:0] verilogPut_KeyCompares_2_429;
  reg [3-1:0] verilogPut_KeyCollapse_2_430;
  reg [64-1:0] verilogPut_Data_2_431;
  reg [64-1:0] verilogPut_Key_3_432;
  reg [1-1:0] verilogPut_KeyCompares_3_433;
  reg [3-1:0] verilogPut_KeyCollapse_3_434;
  reg [64-1:0] verilogPut_Data_3_435;
  reg [1-1:0] verilogPut_Found_436;
  reg [64-1:0] verilogPut_Key_437;
  reg [64-1:0] verilogPut_FoundKey_438;
  reg [64-1:0] verilogPut_Data_439;
  reg [4-1:0] verilogPut_BtreeIndex_440;
  reg [3-1:0] verilogPut_StuckIndex_441;
  reg [1-1:0] verilogPut_MergeSuccess_442;
  reg [4-1:0] verilogPut_index_443;
  reg [3-1:0] verilogPut_size_444;
  reg [1-1:0] verilogPut_isLeaf_445;
  reg [4-1:0] verilogPut_nextFree_446;
  reg [64-1:0] verilogPut_Key_0_447;
  reg [1-1:0] verilogPut_KeyCompares_0_448;
  reg [3-1:0] verilogPut_KeyCollapse_0_449;
  reg [64-1:0] verilogPut_Data_0_450;
  reg [64-1:0] verilogPut_Key_1_451;
  reg [1-1:0] verilogPut_KeyCompares_1_452;
  reg [3-1:0] verilogPut_KeyCollapse_1_453;
  reg [64-1:0] verilogPut_Data_1_454;
  reg [64-1:0] verilogPut_Key_2_455;
  reg [1-1:0] verilogPut_KeyCompares_2_456;
  reg [3-1:0] verilogPut_KeyCollapse_2_457;
  reg [64-1:0] verilogPut_Data_2_458;
  reg [64-1:0] verilogPut_Key_3_459;
  reg [1-1:0] verilogPut_KeyCompares_3_460;
  reg [3-1:0] verilogPut_KeyCollapse_3_461;
  reg [64-1:0] verilogPut_Data_3_462;
  reg [1-1:0] verilogPut_Found_463;
  reg [64-1:0] verilogPut_Key_464;
  reg [64-1:0] verilogPut_FoundKey_465;
  reg [64-1:0] verilogPut_Data_466;
  reg [4-1:0] verilogPut_BtreeIndex_467;
  reg [3-1:0] verilogPut_StuckIndex_468;
  reg [1-1:0] verilogPut_MergeSuccess_469;
  reg [4-1:0] verilogPut_index_470;
  reg [3-1:0] verilogPut_size_471;
  reg [1-1:0] verilogPut_isLeaf_472;
  reg [4-1:0] verilogPut_nextFree_473;
  reg [64-1:0] verilogPut_Key_0_474;
  reg [1-1:0] verilogPut_KeyCompares_0_475;
  reg [3-1:0] verilogPut_KeyCollapse_0_476;
  reg [64-1:0] verilogPut_Data_0_477;
  reg [64-1:0] verilogPut_Key_1_478;
  reg [1-1:0] verilogPut_KeyCompares_1_479;
  reg [3-1:0] verilogPut_KeyCollapse_1_480;
  reg [64-1:0] verilogPut_Data_1_481;
  reg [64-1:0] verilogPut_Key_2_482;
  reg [1-1:0] verilogPut_KeyCompares_2_483;
  reg [3-1:0] verilogPut_KeyCollapse_2_484;
  reg [64-1:0] verilogPut_Data_2_485;
  reg [64-1:0] verilogPut_Key_3_486;
  reg [1-1:0] verilogPut_KeyCompares_3_487;
  reg [3-1:0] verilogPut_KeyCollapse_3_488;
  reg [64-1:0] verilogPut_Data_3_489;
  reg [1-1:0] verilogPut_Found_490;
  reg [64-1:0] verilogPut_Key_491;
  reg [64-1:0] verilogPut_FoundKey_492;
  reg [64-1:0] verilogPut_Data_493;
  reg [4-1:0] verilogPut_BtreeIndex_494;
  reg [3-1:0] verilogPut_StuckIndex_495;
  reg [1-1:0] verilogPut_MergeSuccess_496;
  reg [4-1:0] verilogPut_childIndex_497;
  reg [4-1:0] verilogPut_leftIndex_498;
  reg [64-1:0] verilogPut_midKey_499;
  reg [4-1:0] verilogPut_root_500;
  reg [4-1:0] verilogPut_next_501;
  reg [1-1:0] verilogPut_isLeaf_502;
  reg [1-1:0] verilogPut_isFree_503;
  reg [3-1:0] verilogPut_i_504;
  reg [1-1:0] verilogPut_notFull_505;
  reg [4-1:0] verilogPut_index_506;
  reg [3-1:0] verilogPut_size_507;
  reg [1-1:0] verilogPut_isLeaf_508;
  reg [4-1:0] verilogPut_nextFree_509;
  reg [64-1:0] verilogPut_Key_0_510;
  reg [1-1:0] verilogPut_KeyCompares_0_511;
  reg [3-1:0] verilogPut_KeyCollapse_0_512;
  reg [64-1:0] verilogPut_Data_0_513;
  reg [64-1:0] verilogPut_Key_1_514;
  reg [1-1:0] verilogPut_KeyCompares_1_515;
  reg [3-1:0] verilogPut_KeyCollapse_1_516;
  reg [64-1:0] verilogPut_Data_1_517;
  reg [64-1:0] verilogPut_Key_2_518;
  reg [1-1:0] verilogPut_KeyCompares_2_519;
  reg [3-1:0] verilogPut_KeyCollapse_2_520;
  reg [64-1:0] verilogPut_Data_2_521;
  reg [64-1:0] verilogPut_Key_3_522;
  reg [1-1:0] verilogPut_KeyCompares_3_523;
  reg [3-1:0] verilogPut_KeyCollapse_3_524;
  reg [64-1:0] verilogPut_Data_3_525;
  reg [1-1:0] verilogPut_Found_526;
  reg [64-1:0] verilogPut_Key_527;
  reg [64-1:0] verilogPut_FoundKey_528;
  reg [64-1:0] verilogPut_Data_529;
  reg [4-1:0] verilogPut_BtreeIndex_530;
  reg [3-1:0] verilogPut_StuckIndex_531;
  reg [1-1:0] verilogPut_MergeSuccess_532;
  reg [4-1:0] verilogPut_index_533;
  reg [3-1:0] verilogPut_size_534;
  reg [1-1:0] verilogPut_isLeaf_535;
  reg [4-1:0] verilogPut_nextFree_536;
  reg [64-1:0] verilogPut_Key_0_537;
  reg [1-1:0] verilogPut_KeyCompares_0_538;
  reg [3-1:0] verilogPut_KeyCollapse_0_539;
  reg [64-1:0] verilogPut_Data_0_540;
  reg [64-1:0] verilogPut_Key_1_541;
  reg [1-1:0] verilogPut_KeyCompares_1_542;
  reg [3-1:0] verilogPut_KeyCollapse_1_543;
  reg [64-1:0] verilogPut_Data_1_544;
  reg [64-1:0] verilogPut_Key_2_545;
  reg [1-1:0] verilogPut_KeyCompares_2_546;
  reg [3-1:0] verilogPut_KeyCollapse_2_547;
  reg [64-1:0] verilogPut_Data_2_548;
  reg [64-1:0] verilogPut_Key_3_549;
  reg [1-1:0] verilogPut_KeyCompares_3_550;
  reg [3-1:0] verilogPut_KeyCollapse_3_551;
  reg [64-1:0] verilogPut_Data_3_552;
  reg [1-1:0] verilogPut_Found_553;
  reg [64-1:0] verilogPut_Key_554;
  reg [64-1:0] verilogPut_FoundKey_555;
  reg [64-1:0] verilogPut_Data_556;
  reg [4-1:0] verilogPut_BtreeIndex_557;
  reg [3-1:0] verilogPut_StuckIndex_558;
  reg [1-1:0] verilogPut_MergeSuccess_559;
  reg [4-1:0] verilogPut_index_560;
  reg [3-1:0] verilogPut_size_561;
  reg [1-1:0] verilogPut_isLeaf_562;
  reg [4-1:0] verilogPut_nextFree_563;
  reg [64-1:0] verilogPut_Key_0_564;
  reg [1-1:0] verilogPut_KeyCompares_0_565;
  reg [3-1:0] verilogPut_KeyCollapse_0_566;
  reg [64-1:0] verilogPut_Data_0_567;
  reg [64-1:0] verilogPut_Key_1_568;
  reg [1-1:0] verilogPut_KeyCompares_1_569;
  reg [3-1:0] verilogPut_KeyCollapse_1_570;
  reg [64-1:0] verilogPut_Data_1_571;
  reg [64-1:0] verilogPut_Key_2_572;
  reg [1-1:0] verilogPut_KeyCompares_2_573;
  reg [3-1:0] verilogPut_KeyCollapse_2_574;
  reg [64-1:0] verilogPut_Data_2_575;
  reg [64-1:0] verilogPut_Key_3_576;
  reg [1-1:0] verilogPut_KeyCompares_3_577;
  reg [3-1:0] verilogPut_KeyCollapse_3_578;
  reg [64-1:0] verilogPut_Data_3_579;
  reg [1-1:0] verilogPut_Found_580;
  reg [64-1:0] verilogPut_Key_581;
  reg [64-1:0] verilogPut_FoundKey_582;
  reg [64-1:0] verilogPut_Data_583;
  reg [4-1:0] verilogPut_BtreeIndex_584;
  reg [3-1:0] verilogPut_StuckIndex_585;
  reg [1-1:0] verilogPut_MergeSuccess_586;
  reg [4-1:0] verilogPut_index_587;
  reg [3-1:0] verilogPut_size_588;
  reg [1-1:0] verilogPut_isLeaf_589;
  reg [4-1:0] verilogPut_nextFree_590;
  reg [64-1:0] verilogPut_Key_0_591;
  reg [1-1:0] verilogPut_KeyCompares_0_592;
  reg [3-1:0] verilogPut_KeyCollapse_0_593;
  reg [64-1:0] verilogPut_Data_0_594;
  reg [64-1:0] verilogPut_Key_1_595;
  reg [1-1:0] verilogPut_KeyCompares_1_596;
  reg [3-1:0] verilogPut_KeyCollapse_1_597;
  reg [64-1:0] verilogPut_Data_1_598;
  reg [64-1:0] verilogPut_Key_2_599;
  reg [1-1:0] verilogPut_KeyCompares_2_600;
  reg [3-1:0] verilogPut_KeyCollapse_2_601;
  reg [64-1:0] verilogPut_Data_2_602;
  reg [64-1:0] verilogPut_Key_3_603;
  reg [1-1:0] verilogPut_KeyCompares_3_604;
  reg [3-1:0] verilogPut_KeyCollapse_3_605;
  reg [64-1:0] verilogPut_Data_3_606;
  reg [1-1:0] verilogPut_Found_607;
  reg [64-1:0] verilogPut_Key_608;
  reg [64-1:0] verilogPut_FoundKey_609;
  reg [64-1:0] verilogPut_Data_610;
  reg [4-1:0] verilogPut_BtreeIndex_611;
  reg [3-1:0] verilogPut_StuckIndex_612;
  reg [1-1:0] verilogPut_MergeSuccess_613;
  reg [64-1:0] verilogPut_childKey_614;
  reg [4-1:0] verilogPut_childData_615;
  reg [4-1:0] verilogPut_indexLeft_616;
  reg [4-1:0] verilogPut_indexRight_617;
  reg [64-1:0] verilogPut_midKey_618;
  reg [4-1:0] verilogPut_root_619;
  reg [4-1:0] verilogPut_next_620;
  reg [1-1:0] verilogPut_isLeaf_621;
  reg [1-1:0] verilogPut_isFree_622;
  reg [4-1:0] verilogPut_index_623;
  reg [3-1:0] verilogPut_size_624;
  reg [1-1:0] verilogPut_isLeaf_625;
  reg [4-1:0] verilogPut_nextFree_626;
  reg [64-1:0] verilogPut_Key_0_627;
  reg [1-1:0] verilogPut_KeyCompares_0_628;
  reg [3-1:0] verilogPut_KeyCollapse_0_629;
  reg [64-1:0] verilogPut_Data_0_630;
  reg [64-1:0] verilogPut_Key_1_631;
  reg [1-1:0] verilogPut_KeyCompares_1_632;
  reg [3-1:0] verilogPut_KeyCollapse_1_633;
  reg [64-1:0] verilogPut_Data_1_634;
  reg [64-1:0] verilogPut_Key_2_635;
  reg [1-1:0] verilogPut_KeyCompares_2_636;
  reg [3-1:0] verilogPut_KeyCollapse_2_637;
  reg [64-1:0] verilogPut_Data_2_638;
  reg [64-1:0] verilogPut_Key_3_639;
  reg [1-1:0] verilogPut_KeyCompares_3_640;
  reg [3-1:0] verilogPut_KeyCollapse_3_641;
  reg [64-1:0] verilogPut_Data_3_642;
  reg [1-1:0] verilogPut_Found_643;
  reg [64-1:0] verilogPut_Key_644;
  reg [64-1:0] verilogPut_FoundKey_645;
  reg [64-1:0] verilogPut_Data_646;
  reg [4-1:0] verilogPut_BtreeIndex_647;
  reg [3-1:0] verilogPut_StuckIndex_648;
  reg [1-1:0] verilogPut_MergeSuccess_649;
  reg [4-1:0] verilogPut_index_650;
  reg [3-1:0] verilogPut_size_651;
  reg [1-1:0] verilogPut_isLeaf_652;
  reg [4-1:0] verilogPut_nextFree_653;
  reg [64-1:0] verilogPut_Key_0_654;
  reg [1-1:0] verilogPut_KeyCompares_0_655;
  reg [3-1:0] verilogPut_KeyCollapse_0_656;
  reg [64-1:0] verilogPut_Data_0_657;
  reg [64-1:0] verilogPut_Key_1_658;
  reg [1-1:0] verilogPut_KeyCompares_1_659;
  reg [3-1:0] verilogPut_KeyCollapse_1_660;
  reg [64-1:0] verilogPut_Data_1_661;
  reg [64-1:0] verilogPut_Key_2_662;
  reg [1-1:0] verilogPut_KeyCompares_2_663;
  reg [3-1:0] verilogPut_KeyCollapse_2_664;
  reg [64-1:0] verilogPut_Data_2_665;
  reg [64-1:0] verilogPut_Key_3_666;
  reg [1-1:0] verilogPut_KeyCompares_3_667;
  reg [3-1:0] verilogPut_KeyCollapse_3_668;
  reg [64-1:0] verilogPut_Data_3_669;
  reg [1-1:0] verilogPut_Found_670;
  reg [64-1:0] verilogPut_Key_671;
  reg [64-1:0] verilogPut_FoundKey_672;
  reg [64-1:0] verilogPut_Data_673;
  reg [4-1:0] verilogPut_BtreeIndex_674;
  reg [3-1:0] verilogPut_StuckIndex_675;
  reg [1-1:0] verilogPut_MergeSuccess_676;
  reg [4-1:0] verilogPut_index_677;
  reg [3-1:0] verilogPut_size_678;
  reg [1-1:0] verilogPut_isLeaf_679;
  reg [4-1:0] verilogPut_nextFree_680;
  reg [64-1:0] verilogPut_Key_0_681;
  reg [1-1:0] verilogPut_KeyCompares_0_682;
  reg [3-1:0] verilogPut_KeyCollapse_0_683;
  reg [64-1:0] verilogPut_Data_0_684;
  reg [64-1:0] verilogPut_Key_1_685;
  reg [1-1:0] verilogPut_KeyCompares_1_686;
  reg [3-1:0] verilogPut_KeyCollapse_1_687;
  reg [64-1:0] verilogPut_Data_1_688;
  reg [64-1:0] verilogPut_Key_2_689;
  reg [1-1:0] verilogPut_KeyCompares_2_690;
  reg [3-1:0] verilogPut_KeyCollapse_2_691;
  reg [64-1:0] verilogPut_Data_2_692;
  reg [64-1:0] verilogPut_Key_3_693;
  reg [1-1:0] verilogPut_KeyCompares_3_694;
  reg [3-1:0] verilogPut_KeyCollapse_3_695;
  reg [64-1:0] verilogPut_Data_3_696;
  reg [1-1:0] verilogPut_Found_697;
  reg [64-1:0] verilogPut_Key_698;
  reg [64-1:0] verilogPut_FoundKey_699;
  reg [64-1:0] verilogPut_Data_700;
  reg [4-1:0] verilogPut_BtreeIndex_701;
  reg [3-1:0] verilogPut_StuckIndex_702;
  reg [1-1:0] verilogPut_MergeSuccess_703;
  reg [4-1:0] verilogPut_index_704;
  reg [3-1:0] verilogPut_size_705;
  reg [1-1:0] verilogPut_isLeaf_706;
  reg [4-1:0] verilogPut_nextFree_707;
  reg [64-1:0] verilogPut_Key_0_708;
  reg [1-1:0] verilogPut_KeyCompares_0_709;
  reg [3-1:0] verilogPut_KeyCollapse_0_710;
  reg [64-1:0] verilogPut_Data_0_711;
  reg [64-1:0] verilogPut_Key_1_712;
  reg [1-1:0] verilogPut_KeyCompares_1_713;
  reg [3-1:0] verilogPut_KeyCollapse_1_714;
  reg [64-1:0] verilogPut_Data_1_715;
  reg [64-1:0] verilogPut_Key_2_716;
  reg [1-1:0] verilogPut_KeyCompares_2_717;
  reg [3-1:0] verilogPut_KeyCollapse_2_718;
  reg [64-1:0] verilogPut_Data_2_719;
  reg [64-1:0] verilogPut_Key_3_720;
  reg [1-1:0] verilogPut_KeyCompares_3_721;
  reg [3-1:0] verilogPut_KeyCollapse_3_722;
  reg [64-1:0] verilogPut_Data_3_723;
  reg [1-1:0] verilogPut_Found_724;
  reg [64-1:0] verilogPut_Key_725;
  reg [64-1:0] verilogPut_FoundKey_726;
  reg [64-1:0] verilogPut_Data_727;
  reg [4-1:0] verilogPut_BtreeIndex_728;
  reg [3-1:0] verilogPut_StuckIndex_729;
  reg [1-1:0] verilogPut_MergeSuccess_730;
  reg [64-1:0] verilogPut_childKey_731;
  reg [4-1:0] verilogPut_childData_732;
  reg [4-1:0] verilogPut_indexLeft_733;
  reg [4-1:0] verilogPut_indexRight_734;
  reg [64-1:0] verilogPut_midKey_735;
  reg [4-1:0] verilogPut_root_736;
  reg [4-1:0] verilogPut_next_737;
  reg [1-1:0] verilogPut_isLeaf_738;
  reg [1-1:0] verilogPut_isFree_739;
  reg [4-1:0] verilogPut_index_740;
  reg [3-1:0] verilogPut_size_741;
  reg [1-1:0] verilogPut_isLeaf_742;
  reg [4-1:0] verilogPut_nextFree_743;
  reg [64-1:0] verilogPut_Key_0_744;
  reg [1-1:0] verilogPut_KeyCompares_0_745;
  reg [3-1:0] verilogPut_KeyCollapse_0_746;
  reg [64-1:0] verilogPut_Data_0_747;
  reg [64-1:0] verilogPut_Key_1_748;
  reg [1-1:0] verilogPut_KeyCompares_1_749;
  reg [3-1:0] verilogPut_KeyCollapse_1_750;
  reg [64-1:0] verilogPut_Data_1_751;
  reg [64-1:0] verilogPut_Key_2_752;
  reg [1-1:0] verilogPut_KeyCompares_2_753;
  reg [3-1:0] verilogPut_KeyCollapse_2_754;
  reg [64-1:0] verilogPut_Data_2_755;
  reg [64-1:0] verilogPut_Key_3_756;
  reg [1-1:0] verilogPut_KeyCompares_3_757;
  reg [3-1:0] verilogPut_KeyCollapse_3_758;
  reg [64-1:0] verilogPut_Data_3_759;
  reg [1-1:0] verilogPut_Found_760;
  reg [64-1:0] verilogPut_Key_761;
  reg [64-1:0] verilogPut_FoundKey_762;
  reg [64-1:0] verilogPut_Data_763;
  reg [4-1:0] verilogPut_BtreeIndex_764;
  reg [3-1:0] verilogPut_StuckIndex_765;
  reg [1-1:0] verilogPut_MergeSuccess_766;
  reg [4-1:0] verilogPut_position_767;
  reg [3-1:0] verilogPut_index_768;
  reg [1-1:0] verilogPut_within_769;
  reg [1-1:0] verilogPut_isLeaf_770;
  reg [4-1:0] verilogPut_index_771;
  reg [3-1:0] verilogPut_size_772;
  reg [1-1:0] verilogPut_isLeaf_773;
  reg [4-1:0] verilogPut_nextFree_774;
  reg [64-1:0] verilogPut_Key_0_775;
  reg [1-1:0] verilogPut_KeyCompares_0_776;
  reg [3-1:0] verilogPut_KeyCollapse_0_777;
  reg [64-1:0] verilogPut_Data_0_778;
  reg [64-1:0] verilogPut_Key_1_779;
  reg [1-1:0] verilogPut_KeyCompares_1_780;
  reg [3-1:0] verilogPut_KeyCollapse_1_781;
  reg [64-1:0] verilogPut_Data_1_782;
  reg [64-1:0] verilogPut_Key_2_783;
  reg [1-1:0] verilogPut_KeyCompares_2_784;
  reg [3-1:0] verilogPut_KeyCollapse_2_785;
  reg [64-1:0] verilogPut_Data_2_786;
  reg [64-1:0] verilogPut_Key_3_787;
  reg [1-1:0] verilogPut_KeyCompares_3_788;
  reg [3-1:0] verilogPut_KeyCollapse_3_789;
  reg [64-1:0] verilogPut_Data_3_790;
  reg [1-1:0] verilogPut_Found_791;
  reg [64-1:0] verilogPut_Key_792;
  reg [64-1:0] verilogPut_FoundKey_793;
  reg [64-1:0] verilogPut_Data_794;
  reg [4-1:0] verilogPut_BtreeIndex_795;
  reg [3-1:0] verilogPut_StuckIndex_796;
  reg [1-1:0] verilogPut_MergeSuccess_797;
  reg [4-1:0] verilogPut_index_798;
  reg [3-1:0] verilogPut_size_799;
  reg [1-1:0] verilogPut_isLeaf_800;
  reg [4-1:0] verilogPut_nextFree_801;
  reg [64-1:0] verilogPut_Key_0_802;
  reg [1-1:0] verilogPut_KeyCompares_0_803;
  reg [3-1:0] verilogPut_KeyCollapse_0_804;
  reg [64-1:0] verilogPut_Data_0_805;
  reg [64-1:0] verilogPut_Key_1_806;
  reg [1-1:0] verilogPut_KeyCompares_1_807;
  reg [3-1:0] verilogPut_KeyCollapse_1_808;
  reg [64-1:0] verilogPut_Data_1_809;
  reg [64-1:0] verilogPut_Key_2_810;
  reg [1-1:0] verilogPut_KeyCompares_2_811;
  reg [3-1:0] verilogPut_KeyCollapse_2_812;
  reg [64-1:0] verilogPut_Data_2_813;
  reg [64-1:0] verilogPut_Key_3_814;
  reg [1-1:0] verilogPut_KeyCompares_3_815;
  reg [3-1:0] verilogPut_KeyCollapse_3_816;
  reg [64-1:0] verilogPut_Data_3_817;
  reg [1-1:0] verilogPut_Found_818;
  reg [64-1:0] verilogPut_Key_819;
  reg [64-1:0] verilogPut_FoundKey_820;
  reg [64-1:0] verilogPut_Data_821;
  reg [4-1:0] verilogPut_BtreeIndex_822;
  reg [3-1:0] verilogPut_StuckIndex_823;
  reg [1-1:0] verilogPut_MergeSuccess_824;
  reg [4-1:0] verilogPut_index_825;
  reg [3-1:0] verilogPut_size_826;
  reg [1-1:0] verilogPut_isLeaf_827;
  reg [4-1:0] verilogPut_nextFree_828;
  reg [64-1:0] verilogPut_Key_0_829;
  reg [1-1:0] verilogPut_KeyCompares_0_830;
  reg [3-1:0] verilogPut_KeyCollapse_0_831;
  reg [64-1:0] verilogPut_Data_0_832;
  reg [64-1:0] verilogPut_Key_1_833;
  reg [1-1:0] verilogPut_KeyCompares_1_834;
  reg [3-1:0] verilogPut_KeyCollapse_1_835;
  reg [64-1:0] verilogPut_Data_1_836;
  reg [64-1:0] verilogPut_Key_2_837;
  reg [1-1:0] verilogPut_KeyCompares_2_838;
  reg [3-1:0] verilogPut_KeyCollapse_2_839;
  reg [64-1:0] verilogPut_Data_2_840;
  reg [64-1:0] verilogPut_Key_3_841;
  reg [1-1:0] verilogPut_KeyCompares_3_842;
  reg [3-1:0] verilogPut_KeyCollapse_3_843;
  reg [64-1:0] verilogPut_Data_3_844;
  reg [1-1:0] verilogPut_Found_845;
  reg [64-1:0] verilogPut_Key_846;
  reg [64-1:0] verilogPut_FoundKey_847;
  reg [64-1:0] verilogPut_Data_848;
  reg [4-1:0] verilogPut_BtreeIndex_849;
  reg [3-1:0] verilogPut_StuckIndex_850;
  reg [1-1:0] verilogPut_MergeSuccess_851;
  reg [64-1:0] verilogPut_childKey_852;
  reg [4-1:0] verilogPut_childData_853;
  reg [4-1:0] verilogPut_indexLeft_854;
  reg [4-1:0] verilogPut_indexRight_855;
  reg [64-1:0] verilogPut_midKey_856;
  reg [1-1:0] verilogPut_success_857;
  reg [1-1:0] verilogPut_test_858;
  reg [4-1:0] verilogPut_next_859;
  reg [4-1:0] verilogPut_root_860;
  reg [1-1:0] verilogPut_isFree_861;
  reg [4-1:0] verilogPut_next_862;
  reg [4-1:0] verilogPut_root_863;
  reg [1-1:0] verilogPut_isFree_864;
  reg [4-1:0] verilogPut_index_865;
  reg [3-1:0] verilogPut_size_866;
  reg [1-1:0] verilogPut_isLeaf_867;
  reg [4-1:0] verilogPut_nextFree_868;
  reg [64-1:0] verilogPut_Key_0_869;
  reg [1-1:0] verilogPut_KeyCompares_0_870;
  reg [3-1:0] verilogPut_KeyCollapse_0_871;
  reg [64-1:0] verilogPut_Data_0_872;
  reg [64-1:0] verilogPut_Key_1_873;
  reg [1-1:0] verilogPut_KeyCompares_1_874;
  reg [3-1:0] verilogPut_KeyCollapse_1_875;
  reg [64-1:0] verilogPut_Data_1_876;
  reg [64-1:0] verilogPut_Key_2_877;
  reg [1-1:0] verilogPut_KeyCompares_2_878;
  reg [3-1:0] verilogPut_KeyCollapse_2_879;
  reg [64-1:0] verilogPut_Data_2_880;
  reg [64-1:0] verilogPut_Key_3_881;
  reg [1-1:0] verilogPut_KeyCompares_3_882;
  reg [3-1:0] verilogPut_KeyCollapse_3_883;
  reg [64-1:0] verilogPut_Data_3_884;
  reg [1-1:0] verilogPut_Found_885;
  reg [64-1:0] verilogPut_Key_886;
  reg [64-1:0] verilogPut_FoundKey_887;
  reg [64-1:0] verilogPut_Data_888;
  reg [4-1:0] verilogPut_BtreeIndex_889;
  reg [3-1:0] verilogPut_StuckIndex_890;
  reg [1-1:0] verilogPut_MergeSuccess_891;
  reg [4-1:0] verilogPut_index_892;
  reg [3-1:0] verilogPut_size_893;
  reg [1-1:0] verilogPut_isLeaf_894;
  reg [4-1:0] verilogPut_nextFree_895;
  reg [64-1:0] verilogPut_Key_0_896;
  reg [1-1:0] verilogPut_KeyCompares_0_897;
  reg [3-1:0] verilogPut_KeyCollapse_0_898;
  reg [64-1:0] verilogPut_Data_0_899;
  reg [64-1:0] verilogPut_Key_1_900;
  reg [1-1:0] verilogPut_KeyCompares_1_901;
  reg [3-1:0] verilogPut_KeyCollapse_1_902;
  reg [64-1:0] verilogPut_Data_1_903;
  reg [64-1:0] verilogPut_Key_2_904;
  reg [1-1:0] verilogPut_KeyCompares_2_905;
  reg [3-1:0] verilogPut_KeyCollapse_2_906;
  reg [64-1:0] verilogPut_Data_2_907;
  reg [64-1:0] verilogPut_Key_3_908;
  reg [1-1:0] verilogPut_KeyCompares_3_909;
  reg [3-1:0] verilogPut_KeyCollapse_3_910;
  reg [64-1:0] verilogPut_Data_3_911;
  reg [1-1:0] verilogPut_Found_912;
  reg [64-1:0] verilogPut_Key_913;
  reg [64-1:0] verilogPut_FoundKey_914;
  reg [64-1:0] verilogPut_Data_915;
  reg [4-1:0] verilogPut_BtreeIndex_916;
  reg [3-1:0] verilogPut_StuckIndex_917;
  reg [1-1:0] verilogPut_MergeSuccess_918;
  reg [4-1:0] verilogPut_index_919;
  reg [3-1:0] verilogPut_size_920;
  reg [1-1:0] verilogPut_isLeaf_921;
  reg [4-1:0] verilogPut_nextFree_922;
  reg [64-1:0] verilogPut_Key_0_923;
  reg [1-1:0] verilogPut_KeyCompares_0_924;
  reg [3-1:0] verilogPut_KeyCollapse_0_925;
  reg [64-1:0] verilogPut_Data_0_926;
  reg [64-1:0] verilogPut_Key_1_927;
  reg [1-1:0] verilogPut_KeyCompares_1_928;
  reg [3-1:0] verilogPut_KeyCollapse_1_929;
  reg [64-1:0] verilogPut_Data_1_930;
  reg [64-1:0] verilogPut_Key_2_931;
  reg [1-1:0] verilogPut_KeyCompares_2_932;
  reg [3-1:0] verilogPut_KeyCollapse_2_933;
  reg [64-1:0] verilogPut_Data_2_934;
  reg [64-1:0] verilogPut_Key_3_935;
  reg [1-1:0] verilogPut_KeyCompares_3_936;
  reg [3-1:0] verilogPut_KeyCollapse_3_937;
  reg [64-1:0] verilogPut_Data_3_938;
  reg [1-1:0] verilogPut_Found_939;
  reg [64-1:0] verilogPut_Key_940;
  reg [64-1:0] verilogPut_FoundKey_941;
  reg [64-1:0] verilogPut_Data_942;
  reg [4-1:0] verilogPut_BtreeIndex_943;
  reg [3-1:0] verilogPut_StuckIndex_944;
  reg [1-1:0] verilogPut_MergeSuccess_945;
  reg [64-1:0] verilogPut_childKey_946;
  reg [3-1:0] verilogPut_leftChild_947;
  reg [3-1:0] verilogPut_rightChild_948;
  reg [4-1:0] verilogPut_childData_949;
  reg [4-1:0] verilogPut_indexLeft_950;
  reg [4-1:0] verilogPut_indexRight_951;
  reg [64-1:0] verilogPut_midKey_952;
  reg [1-1:0] verilogPut_success_953;
  reg [1-1:0] verilogPut_test_954;
  reg [4-1:0] verilogPut_next_955;
  reg [4-1:0] verilogPut_root_956;
  reg [1-1:0] verilogPut_isFree_957;
  reg [4-1:0] verilogPut_next_958;
  reg [4-1:0] verilogPut_root_959;
  reg [1-1:0] verilogPut_isFree_960;
  reg [4-1:0] verilogPut_index_961;
  reg [3-1:0] verilogPut_size_962;
  reg [1-1:0] verilogPut_isLeaf_963;
  reg [4-1:0] verilogPut_nextFree_964;
  reg [64-1:0] verilogPut_Key_0_965;
  reg [1-1:0] verilogPut_KeyCompares_0_966;
  reg [3-1:0] verilogPut_KeyCollapse_0_967;
  reg [64-1:0] verilogPut_Data_0_968;
  reg [64-1:0] verilogPut_Key_1_969;
  reg [1-1:0] verilogPut_KeyCompares_1_970;
  reg [3-1:0] verilogPut_KeyCollapse_1_971;
  reg [64-1:0] verilogPut_Data_1_972;
  reg [64-1:0] verilogPut_Key_2_973;
  reg [1-1:0] verilogPut_KeyCompares_2_974;
  reg [3-1:0] verilogPut_KeyCollapse_2_975;
  reg [64-1:0] verilogPut_Data_2_976;
  reg [64-1:0] verilogPut_Key_3_977;
  reg [1-1:0] verilogPut_KeyCompares_3_978;
  reg [3-1:0] verilogPut_KeyCollapse_3_979;
  reg [64-1:0] verilogPut_Data_3_980;
  reg [1-1:0] verilogPut_Found_981;
  reg [64-1:0] verilogPut_Key_982;
  reg [64-1:0] verilogPut_FoundKey_983;
  reg [64-1:0] verilogPut_Data_984;
  reg [4-1:0] verilogPut_BtreeIndex_985;
  reg [3-1:0] verilogPut_StuckIndex_986;
  reg [1-1:0] verilogPut_MergeSuccess_987;
  reg [4-1:0] verilogPut_index_988;
  reg [3-1:0] verilogPut_size_989;
  reg [1-1:0] verilogPut_isLeaf_990;
  reg [4-1:0] verilogPut_nextFree_991;
  reg [64-1:0] verilogPut_Key_0_992;
  reg [1-1:0] verilogPut_KeyCompares_0_993;
  reg [3-1:0] verilogPut_KeyCollapse_0_994;
  reg [64-1:0] verilogPut_Data_0_995;
  reg [64-1:0] verilogPut_Key_1_996;
  reg [1-1:0] verilogPut_KeyCompares_1_997;
  reg [3-1:0] verilogPut_KeyCollapse_1_998;
  reg [64-1:0] verilogPut_Data_1_999;
  reg [64-1:0] verilogPut_Key_2_1000;
  reg [1-1:0] verilogPut_KeyCompares_2_1001;
  reg [3-1:0] verilogPut_KeyCollapse_2_1002;
  reg [64-1:0] verilogPut_Data_2_1003;
  reg [64-1:0] verilogPut_Key_3_1004;
  reg [1-1:0] verilogPut_KeyCompares_3_1005;
  reg [3-1:0] verilogPut_KeyCollapse_3_1006;
  reg [64-1:0] verilogPut_Data_3_1007;
  reg [1-1:0] verilogPut_Found_1008;
  reg [64-1:0] verilogPut_Key_1009;
  reg [64-1:0] verilogPut_FoundKey_1010;
  reg [64-1:0] verilogPut_Data_1011;
  reg [4-1:0] verilogPut_BtreeIndex_1012;
  reg [3-1:0] verilogPut_StuckIndex_1013;
  reg [1-1:0] verilogPut_MergeSuccess_1014;
  reg [64-1:0] verilogPut_childKey_1015;
  reg [3-1:0] verilogPut_size_1016;
  reg [4-1:0] verilogPut_childData_1017;
  reg [4-1:0] verilogPut_indexLeft_1018;
  reg [4-1:0] verilogPut_indexRight_1019;
  reg [64-1:0] verilogPut_midKey_1020;
  reg [1-1:0] verilogPut_success_1021;
  reg [1-1:0] verilogPut_test_1022;
  reg [4-1:0] verilogPut_next_1023;
  reg [4-1:0] verilogPut_root_1024;
  reg [1-1:0] verilogPut_isFree_1025;
  reg [4-1:0] verilogPut_index_1026;
  reg [3-1:0] verilogPut_size_1027;
  reg [1-1:0] verilogPut_isLeaf_1028;
  reg [4-1:0] verilogPut_nextFree_1029;
  reg [64-1:0] verilogPut_Key_0_1030;
  reg [1-1:0] verilogPut_KeyCompares_0_1031;
  reg [3-1:0] verilogPut_KeyCollapse_0_1032;
  reg [64-1:0] verilogPut_Data_0_1033;
  reg [64-1:0] verilogPut_Key_1_1034;
  reg [1-1:0] verilogPut_KeyCompares_1_1035;
  reg [3-1:0] verilogPut_KeyCollapse_1_1036;
  reg [64-1:0] verilogPut_Data_1_1037;
  reg [64-1:0] verilogPut_Key_2_1038;
  reg [1-1:0] verilogPut_KeyCompares_2_1039;
  reg [3-1:0] verilogPut_KeyCollapse_2_1040;
  reg [64-1:0] verilogPut_Data_2_1041;
  reg [64-1:0] verilogPut_Key_3_1042;
  reg [1-1:0] verilogPut_KeyCompares_3_1043;
  reg [3-1:0] verilogPut_KeyCollapse_3_1044;
  reg [64-1:0] verilogPut_Data_3_1045;
  reg [1-1:0] verilogPut_Found_1046;
  reg [64-1:0] verilogPut_Key_1047;
  reg [64-1:0] verilogPut_FoundKey_1048;
  reg [64-1:0] verilogPut_Data_1049;
  reg [4-1:0] verilogPut_BtreeIndex_1050;
  reg [3-1:0] verilogPut_StuckIndex_1051;
  reg [1-1:0] verilogPut_MergeSuccess_1052;
  reg [4-1:0] verilogPut_index_1053;
  reg [3-1:0] verilogPut_size_1054;
  reg [1-1:0] verilogPut_isLeaf_1055;
  reg [4-1:0] verilogPut_nextFree_1056;
  reg [64-1:0] verilogPut_Key_0_1057;
  reg [1-1:0] verilogPut_KeyCompares_0_1058;
  reg [3-1:0] verilogPut_KeyCollapse_0_1059;
  reg [64-1:0] verilogPut_Data_0_1060;
  reg [64-1:0] verilogPut_Key_1_1061;
  reg [1-1:0] verilogPut_KeyCompares_1_1062;
  reg [3-1:0] verilogPut_KeyCollapse_1_1063;
  reg [64-1:0] verilogPut_Data_1_1064;
  reg [64-1:0] verilogPut_Key_2_1065;
  reg [1-1:0] verilogPut_KeyCompares_2_1066;
  reg [3-1:0] verilogPut_KeyCollapse_2_1067;
  reg [64-1:0] verilogPut_Data_2_1068;
  reg [64-1:0] verilogPut_Key_3_1069;
  reg [1-1:0] verilogPut_KeyCompares_3_1070;
  reg [3-1:0] verilogPut_KeyCollapse_3_1071;
  reg [64-1:0] verilogPut_Data_3_1072;
  reg [1-1:0] verilogPut_Found_1073;
  reg [64-1:0] verilogPut_Key_1074;
  reg [64-1:0] verilogPut_FoundKey_1075;
  reg [64-1:0] verilogPut_Data_1076;
  reg [4-1:0] verilogPut_BtreeIndex_1077;
  reg [3-1:0] verilogPut_StuckIndex_1078;
  reg [1-1:0] verilogPut_MergeSuccess_1079;
  reg [64-1:0] verilogPut_childKey_1080;
  reg [3-1:0] verilogPut_size_1081;
  reg [4-1:0] verilogPut_childData_1082;
  reg [4-1:0] verilogPut_indexLeft_1083;
  reg [4-1:0] verilogPut_indexRight_1084;
  reg [64-1:0] verilogPut_midKey_1085;
  reg [1-1:0] verilogPut_success_1086;
  reg [1-1:0] verilogPut_test_1087;
  reg [4-1:0] verilogPut_next_1088;
  reg [4-1:0] verilogPut_root_1089;
  reg [1-1:0] verilogPut_isFree_1090;
  reg [4-1:0] verilogPut_index_1091;
  reg [3-1:0] verilogPut_size_1092;
  reg [1-1:0] verilogPut_isLeaf_1093;
  reg [4-1:0] verilogPut_nextFree_1094;
  reg [64-1:0] verilogPut_Key_0_1095;
  reg [1-1:0] verilogPut_KeyCompares_0_1096;
  reg [3-1:0] verilogPut_KeyCollapse_0_1097;
  reg [64-1:0] verilogPut_Data_0_1098;
  reg [64-1:0] verilogPut_Key_1_1099;
  reg [1-1:0] verilogPut_KeyCompares_1_1100;
  reg [3-1:0] verilogPut_KeyCollapse_1_1101;
  reg [64-1:0] verilogPut_Data_1_1102;
  reg [64-1:0] verilogPut_Key_2_1103;
  reg [1-1:0] verilogPut_KeyCompares_2_1104;
  reg [3-1:0] verilogPut_KeyCollapse_2_1105;
  reg [64-1:0] verilogPut_Data_2_1106;
  reg [64-1:0] verilogPut_Key_3_1107;
  reg [1-1:0] verilogPut_KeyCompares_3_1108;
  reg [3-1:0] verilogPut_KeyCollapse_3_1109;
  reg [64-1:0] verilogPut_Data_3_1110;
  reg [1-1:0] verilogPut_Found_1111;
  reg [64-1:0] verilogPut_Key_1112;
  reg [64-1:0] verilogPut_FoundKey_1113;
  reg [64-1:0] verilogPut_Data_1114;
  reg [4-1:0] verilogPut_BtreeIndex_1115;
  reg [3-1:0] verilogPut_StuckIndex_1116;
  reg [1-1:0] verilogPut_MergeSuccess_1117;
  reg [4-1:0] verilogPut_index_1118;
  reg [3-1:0] verilogPut_size_1119;
  reg [1-1:0] verilogPut_isLeaf_1120;
  reg [4-1:0] verilogPut_nextFree_1121;
  reg [64-1:0] verilogPut_Key_0_1122;
  reg [1-1:0] verilogPut_KeyCompares_0_1123;
  reg [3-1:0] verilogPut_KeyCollapse_0_1124;
  reg [64-1:0] verilogPut_Data_0_1125;
  reg [64-1:0] verilogPut_Key_1_1126;
  reg [1-1:0] verilogPut_KeyCompares_1_1127;
  reg [3-1:0] verilogPut_KeyCollapse_1_1128;
  reg [64-1:0] verilogPut_Data_1_1129;
  reg [64-1:0] verilogPut_Key_2_1130;
  reg [1-1:0] verilogPut_KeyCompares_2_1131;
  reg [3-1:0] verilogPut_KeyCollapse_2_1132;
  reg [64-1:0] verilogPut_Data_2_1133;
  reg [64-1:0] verilogPut_Key_3_1134;
  reg [1-1:0] verilogPut_KeyCompares_3_1135;
  reg [3-1:0] verilogPut_KeyCollapse_3_1136;
  reg [64-1:0] verilogPut_Data_3_1137;
  reg [1-1:0] verilogPut_Found_1138;
  reg [64-1:0] verilogPut_Key_1139;
  reg [64-1:0] verilogPut_FoundKey_1140;
  reg [64-1:0] verilogPut_Data_1141;
  reg [4-1:0] verilogPut_BtreeIndex_1142;
  reg [3-1:0] verilogPut_StuckIndex_1143;
  reg [1-1:0] verilogPut_MergeSuccess_1144;
  reg [64-1:0] verilogPut_childKey_1145;
  reg [4-1:0] verilogPut_childData_1146;
  reg [4-1:0] verilogPut_indexLeft_1147;
  reg [4-1:0] verilogPut_indexRight_1148;
  reg [64-1:0] verilogPut_midKey_1149;
  reg [1-1:0] verilogPut_success_1150;
  reg [1-1:0] verilogPut_test_1151;
  reg [4-1:0] verilogPut_next_1152;
  reg [4-1:0] verilogPut_root_1153;
  reg [1-1:0] verilogPut_isFree_1154;
  reg [4-1:0] verilogPut_index_1155;
  reg [3-1:0] verilogPut_size_1156;
  reg [1-1:0] verilogPut_isLeaf_1157;
  reg [4-1:0] verilogPut_nextFree_1158;
  reg [64-1:0] verilogPut_Key_0_1159;
  reg [1-1:0] verilogPut_KeyCompares_0_1160;
  reg [3-1:0] verilogPut_KeyCollapse_0_1161;
  reg [64-1:0] verilogPut_Data_0_1162;
  reg [64-1:0] verilogPut_Key_1_1163;
  reg [1-1:0] verilogPut_KeyCompares_1_1164;
  reg [3-1:0] verilogPut_KeyCollapse_1_1165;
  reg [64-1:0] verilogPut_Data_1_1166;
  reg [64-1:0] verilogPut_Key_2_1167;
  reg [1-1:0] verilogPut_KeyCompares_2_1168;
  reg [3-1:0] verilogPut_KeyCollapse_2_1169;
  reg [64-1:0] verilogPut_Data_2_1170;
  reg [64-1:0] verilogPut_Key_3_1171;
  reg [1-1:0] verilogPut_KeyCompares_3_1172;
  reg [3-1:0] verilogPut_KeyCollapse_3_1173;
  reg [64-1:0] verilogPut_Data_3_1174;
  reg [1-1:0] verilogPut_Found_1175;
  reg [64-1:0] verilogPut_Key_1176;
  reg [64-1:0] verilogPut_FoundKey_1177;
  reg [64-1:0] verilogPut_Data_1178;
  reg [4-1:0] verilogPut_BtreeIndex_1179;
  reg [3-1:0] verilogPut_StuckIndex_1180;
  reg [1-1:0] verilogPut_MergeSuccess_1181;
  reg [4-1:0] verilogPut_index_1182;
  reg [3-1:0] verilogPut_size_1183;
  reg [1-1:0] verilogPut_isLeaf_1184;
  reg [4-1:0] verilogPut_nextFree_1185;
  reg [64-1:0] verilogPut_Key_0_1186;
  reg [1-1:0] verilogPut_KeyCompares_0_1187;
  reg [3-1:0] verilogPut_KeyCollapse_0_1188;
  reg [64-1:0] verilogPut_Data_0_1189;
  reg [64-1:0] verilogPut_Key_1_1190;
  reg [1-1:0] verilogPut_KeyCompares_1_1191;
  reg [3-1:0] verilogPut_KeyCollapse_1_1192;
  reg [64-1:0] verilogPut_Data_1_1193;
  reg [64-1:0] verilogPut_Key_2_1194;
  reg [1-1:0] verilogPut_KeyCompares_2_1195;
  reg [3-1:0] verilogPut_KeyCollapse_2_1196;
  reg [64-1:0] verilogPut_Data_2_1197;
  reg [64-1:0] verilogPut_Key_3_1198;
  reg [1-1:0] verilogPut_KeyCompares_3_1199;
  reg [3-1:0] verilogPut_KeyCollapse_3_1200;
  reg [64-1:0] verilogPut_Data_3_1201;
  reg [1-1:0] verilogPut_Found_1202;
  reg [64-1:0] verilogPut_Key_1203;
  reg [64-1:0] verilogPut_FoundKey_1204;
  reg [64-1:0] verilogPut_Data_1205;
  reg [4-1:0] verilogPut_BtreeIndex_1206;
  reg [3-1:0] verilogPut_StuckIndex_1207;
  reg [1-1:0] verilogPut_MergeSuccess_1208;
  reg [64-1:0] verilogPut_childKey_1209;
  reg [3-1:0] verilogPut_leftChild_1210;
  reg [3-1:0] verilogPut_rightChild_1211;
  reg [4-1:0] verilogPut_childData_1212;
  reg [4-1:0] verilogPut_indexLeft_1213;
  reg [4-1:0] verilogPut_indexRight_1214;
  reg [64-1:0] verilogPut_midKey_1215;
  reg [1-1:0] verilogPut_success_1216;
  reg [1-1:0] verilogPut_test_1217;
  reg [4-1:0] verilogPut_next_1218;
  reg [4-1:0] verilogPut_root_1219;
  reg [1-1:0] verilogPut_isFree_1220;
  reg [4-1:0] verilogPut_index_1221;
  reg [3-1:0] verilogPut_size_1222;
  reg [1-1:0] verilogPut_isLeaf_1223;
  reg [4-1:0] verilogPut_nextFree_1224;
  reg [64-1:0] verilogPut_Key_0_1225;
  reg [1-1:0] verilogPut_KeyCompares_0_1226;
  reg [3-1:0] verilogPut_KeyCollapse_0_1227;
  reg [64-1:0] verilogPut_Data_0_1228;
  reg [64-1:0] verilogPut_Key_1_1229;
  reg [1-1:0] verilogPut_KeyCompares_1_1230;
  reg [3-1:0] verilogPut_KeyCollapse_1_1231;
  reg [64-1:0] verilogPut_Data_1_1232;
  reg [64-1:0] verilogPut_Key_2_1233;
  reg [1-1:0] verilogPut_KeyCompares_2_1234;
  reg [3-1:0] verilogPut_KeyCollapse_2_1235;
  reg [64-1:0] verilogPut_Data_2_1236;
  reg [64-1:0] verilogPut_Key_3_1237;
  reg [1-1:0] verilogPut_KeyCompares_3_1238;
  reg [3-1:0] verilogPut_KeyCollapse_3_1239;
  reg [64-1:0] verilogPut_Data_3_1240;
  reg [1-1:0] verilogPut_Found_1241;
  reg [64-1:0] verilogPut_Key_1242;
  reg [64-1:0] verilogPut_FoundKey_1243;
  reg [64-1:0] verilogPut_Data_1244;
  reg [4-1:0] verilogPut_BtreeIndex_1245;
  reg [3-1:0] verilogPut_StuckIndex_1246;
  reg [1-1:0] verilogPut_MergeSuccess_1247;
  reg [4-1:0] verilogPut_index_1248;
  reg [3-1:0] verilogPut_size_1249;
  reg [1-1:0] verilogPut_isLeaf_1250;
  reg [4-1:0] verilogPut_nextFree_1251;
  reg [64-1:0] verilogPut_Key_0_1252;
  reg [1-1:0] verilogPut_KeyCompares_0_1253;
  reg [3-1:0] verilogPut_KeyCollapse_0_1254;
  reg [64-1:0] verilogPut_Data_0_1255;
  reg [64-1:0] verilogPut_Key_1_1256;
  reg [1-1:0] verilogPut_KeyCompares_1_1257;
  reg [3-1:0] verilogPut_KeyCollapse_1_1258;
  reg [64-1:0] verilogPut_Data_1_1259;
  reg [64-1:0] verilogPut_Key_2_1260;
  reg [1-1:0] verilogPut_KeyCompares_2_1261;
  reg [3-1:0] verilogPut_KeyCollapse_2_1262;
  reg [64-1:0] verilogPut_Data_2_1263;
  reg [64-1:0] verilogPut_Key_3_1264;
  reg [1-1:0] verilogPut_KeyCompares_3_1265;
  reg [3-1:0] verilogPut_KeyCollapse_3_1266;
  reg [64-1:0] verilogPut_Data_3_1267;
  reg [1-1:0] verilogPut_Found_1268;
  reg [64-1:0] verilogPut_Key_1269;
  reg [64-1:0] verilogPut_FoundKey_1270;
  reg [64-1:0] verilogPut_Data_1271;
  reg [4-1:0] verilogPut_BtreeIndex_1272;
  reg [3-1:0] verilogPut_StuckIndex_1273;
  reg [1-1:0] verilogPut_MergeSuccess_1274;
  reg [64-1:0] verilogPut_childKey_1275;
  reg [4-1:0] verilogPut_childData_1276;
  reg [4-1:0] verilogPut_indexLeft_1277;
  reg [4-1:0] verilogPut_indexRight_1278;
  reg [64-1:0] verilogPut_midKey_1279;
  reg [1-1:0] verilogPut_success_1280;
  reg [1-1:0] verilogPut_test_1281;
  reg [4-1:0] verilogPut_next_1282;
  reg [4-1:0] verilogPut_root_1283;
  reg [1-1:0] verilogPut_isFree_1284;
  reg [4-1:0] verilogPut_index_1285;
  reg [3-1:0] verilogPut_size_1286;
  reg [1-1:0] verilogPut_isLeaf_1287;
  reg [4-1:0] verilogPut_nextFree_1288;
  reg [64-1:0] verilogPut_Key_0_1289;
  reg [1-1:0] verilogPut_KeyCompares_0_1290;
  reg [3-1:0] verilogPut_KeyCollapse_0_1291;
  reg [64-1:0] verilogPut_Data_0_1292;
  reg [64-1:0] verilogPut_Key_1_1293;
  reg [1-1:0] verilogPut_KeyCompares_1_1294;
  reg [3-1:0] verilogPut_KeyCollapse_1_1295;
  reg [64-1:0] verilogPut_Data_1_1296;
  reg [64-1:0] verilogPut_Key_2_1297;
  reg [1-1:0] verilogPut_KeyCompares_2_1298;
  reg [3-1:0] verilogPut_KeyCollapse_2_1299;
  reg [64-1:0] verilogPut_Data_2_1300;
  reg [64-1:0] verilogPut_Key_3_1301;
  reg [1-1:0] verilogPut_KeyCompares_3_1302;
  reg [3-1:0] verilogPut_KeyCollapse_3_1303;
  reg [64-1:0] verilogPut_Data_3_1304;
  reg [1-1:0] verilogPut_Found_1305;
  reg [64-1:0] verilogPut_Key_1306;
  reg [64-1:0] verilogPut_FoundKey_1307;
  reg [64-1:0] verilogPut_Data_1308;
  reg [4-1:0] verilogPut_BtreeIndex_1309;
  reg [3-1:0] verilogPut_StuckIndex_1310;
  reg [1-1:0] verilogPut_MergeSuccess_1311;
  reg [4-1:0] verilogPut_index_1312;
  reg [3-1:0] verilogPut_size_1313;
  reg [1-1:0] verilogPut_isLeaf_1314;
  reg [4-1:0] verilogPut_nextFree_1315;
  reg [64-1:0] verilogPut_Key_0_1316;
  reg [1-1:0] verilogPut_KeyCompares_0_1317;
  reg [3-1:0] verilogPut_KeyCollapse_0_1318;
  reg [64-1:0] verilogPut_Data_0_1319;
  reg [64-1:0] verilogPut_Key_1_1320;
  reg [1-1:0] verilogPut_KeyCompares_1_1321;
  reg [3-1:0] verilogPut_KeyCollapse_1_1322;
  reg [64-1:0] verilogPut_Data_1_1323;
  reg [64-1:0] verilogPut_Key_2_1324;
  reg [1-1:0] verilogPut_KeyCompares_2_1325;
  reg [3-1:0] verilogPut_KeyCollapse_2_1326;
  reg [64-1:0] verilogPut_Data_2_1327;
  reg [64-1:0] verilogPut_Key_3_1328;
  reg [1-1:0] verilogPut_KeyCompares_3_1329;
  reg [3-1:0] verilogPut_KeyCollapse_3_1330;
  reg [64-1:0] verilogPut_Data_3_1331;
  reg [1-1:0] verilogPut_Found_1332;
  reg [64-1:0] verilogPut_Key_1333;
  reg [64-1:0] verilogPut_FoundKey_1334;
  reg [64-1:0] verilogPut_Data_1335;
  reg [4-1:0] verilogPut_BtreeIndex_1336;
  reg [3-1:0] verilogPut_StuckIndex_1337;
  reg [1-1:0] verilogPut_MergeSuccess_1338;
  reg [64-1:0] verilogPut_childKey_1339;
  reg [3-1:0] verilogPut_leftChild_1340;
  reg [3-1:0] verilogPut_rightChild_1341;
  reg [4-1:0] verilogPut_childData_1342;
  reg [4-1:0] verilogPut_indexLeft_1343;
  reg [4-1:0] verilogPut_indexRight_1344;
  reg [64-1:0] verilogPut_midKey_1345;
  reg [1-1:0] verilogPut_success_1346;
  reg [1-1:0] verilogPut_test_1347;
  reg [4-1:0] verilogPut_next_1348;
  reg [4-1:0] verilogPut_root_1349;
  reg [1-1:0] verilogPut_isFree_1350;
  reg [4-1:0] verilogPut_index_1351;
  reg [3-1:0] verilogPut_size_1352;
  reg [1-1:0] verilogPut_isLeaf_1353;
  reg [4-1:0] verilogPut_nextFree_1354;
  reg [64-1:0] verilogPut_Key_0_1355;
  reg [1-1:0] verilogPut_KeyCompares_0_1356;
  reg [3-1:0] verilogPut_KeyCollapse_0_1357;
  reg [64-1:0] verilogPut_Data_0_1358;
  reg [64-1:0] verilogPut_Key_1_1359;
  reg [1-1:0] verilogPut_KeyCompares_1_1360;
  reg [3-1:0] verilogPut_KeyCollapse_1_1361;
  reg [64-1:0] verilogPut_Data_1_1362;
  reg [64-1:0] verilogPut_Key_2_1363;
  reg [1-1:0] verilogPut_KeyCompares_2_1364;
  reg [3-1:0] verilogPut_KeyCollapse_2_1365;
  reg [64-1:0] verilogPut_Data_2_1366;
  reg [64-1:0] verilogPut_Key_3_1367;
  reg [1-1:0] verilogPut_KeyCompares_3_1368;
  reg [3-1:0] verilogPut_KeyCollapse_3_1369;
  reg [64-1:0] verilogPut_Data_3_1370;
  reg [1-1:0] verilogPut_Found_1371;
  reg [64-1:0] verilogPut_Key_1372;
  reg [64-1:0] verilogPut_FoundKey_1373;
  reg [64-1:0] verilogPut_Data_1374;
  reg [4-1:0] verilogPut_BtreeIndex_1375;
  reg [3-1:0] verilogPut_StuckIndex_1376;
  reg [1-1:0] verilogPut_MergeSuccess_1377;
  reg [4-1:0] verilogPut_index_1378;
  reg [3-1:0] verilogPut_size_1379;
  reg [1-1:0] verilogPut_isLeaf_1380;
  reg [4-1:0] verilogPut_nextFree_1381;
  reg [64-1:0] verilogPut_Key_0_1382;
  reg [1-1:0] verilogPut_KeyCompares_0_1383;
  reg [3-1:0] verilogPut_KeyCollapse_0_1384;
  reg [64-1:0] verilogPut_Data_0_1385;
  reg [64-1:0] verilogPut_Key_1_1386;
  reg [1-1:0] verilogPut_KeyCompares_1_1387;
  reg [3-1:0] verilogPut_KeyCollapse_1_1388;
  reg [64-1:0] verilogPut_Data_1_1389;
  reg [64-1:0] verilogPut_Key_2_1390;
  reg [1-1:0] verilogPut_KeyCompares_2_1391;
  reg [3-1:0] verilogPut_KeyCollapse_2_1392;
  reg [64-1:0] verilogPut_Data_2_1393;
  reg [64-1:0] verilogPut_Key_3_1394;
  reg [1-1:0] verilogPut_KeyCompares_3_1395;
  reg [3-1:0] verilogPut_KeyCollapse_3_1396;
  reg [64-1:0] verilogPut_Data_3_1397;
  reg [1-1:0] verilogPut_Found_1398;
  reg [64-1:0] verilogPut_Key_1399;
  reg [64-1:0] verilogPut_FoundKey_1400;
  reg [64-1:0] verilogPut_Data_1401;
  reg [4-1:0] verilogPut_BtreeIndex_1402;
  reg [3-1:0] verilogPut_StuckIndex_1403;
  reg [1-1:0] verilogPut_MergeSuccess_1404;
  reg [64-1:0] verilogPut_childKey_1405;
  reg [4-1:0] verilogPut_childData_1406;
  reg [4-1:0] verilogPut_indexLeft_1407;
  reg [4-1:0] verilogPut_indexRight_1408;
  reg [64-1:0] verilogPut_midKey_1409;
  reg [1-1:0] verilogPut_success_1410;
  reg [1-1:0] verilogPut_test_1411;
  reg [4-1:0] verilogPut_next_1412;
  reg [4-1:0] verilogPut_root_1413;
  reg [1-1:0] verilogPut_isFree_1414;
  reg [4-1:0] verilogPut_index_1415;
  reg [3-1:0] verilogPut_size_1416;
  reg [1-1:0] verilogPut_isLeaf_1417;
  reg [4-1:0] verilogPut_nextFree_1418;
  reg [64-1:0] verilogPut_Key_0_1419;
  reg [1-1:0] verilogPut_KeyCompares_0_1420;
  reg [3-1:0] verilogPut_KeyCollapse_0_1421;
  reg [64-1:0] verilogPut_Data_0_1422;
  reg [64-1:0] verilogPut_Key_1_1423;
  reg [1-1:0] verilogPut_KeyCompares_1_1424;
  reg [3-1:0] verilogPut_KeyCollapse_1_1425;
  reg [64-1:0] verilogPut_Data_1_1426;
  reg [64-1:0] verilogPut_Key_2_1427;
  reg [1-1:0] verilogPut_KeyCompares_2_1428;
  reg [3-1:0] verilogPut_KeyCollapse_2_1429;
  reg [64-1:0] verilogPut_Data_2_1430;
  reg [64-1:0] verilogPut_Key_3_1431;
  reg [1-1:0] verilogPut_KeyCompares_3_1432;
  reg [3-1:0] verilogPut_KeyCollapse_3_1433;
  reg [64-1:0] verilogPut_Data_3_1434;
  reg [1-1:0] verilogPut_Found_1435;
  reg [64-1:0] verilogPut_Key_1436;
  reg [64-1:0] verilogPut_FoundKey_1437;
  reg [64-1:0] verilogPut_Data_1438;
  reg [4-1:0] verilogPut_BtreeIndex_1439;
  reg [3-1:0] verilogPut_StuckIndex_1440;
  reg [1-1:0] verilogPut_MergeSuccess_1441;
  reg [4-1:0] verilogPut_index_1442;
  reg [3-1:0] verilogPut_size_1443;
  reg [1-1:0] verilogPut_isLeaf_1444;
  reg [4-1:0] verilogPut_nextFree_1445;
  reg [64-1:0] verilogPut_Key_0_1446;
  reg [1-1:0] verilogPut_KeyCompares_0_1447;
  reg [3-1:0] verilogPut_KeyCollapse_0_1448;
  reg [64-1:0] verilogPut_Data_0_1449;
  reg [64-1:0] verilogPut_Key_1_1450;
  reg [1-1:0] verilogPut_KeyCompares_1_1451;
  reg [3-1:0] verilogPut_KeyCollapse_1_1452;
  reg [64-1:0] verilogPut_Data_1_1453;
  reg [64-1:0] verilogPut_Key_2_1454;
  reg [1-1:0] verilogPut_KeyCompares_2_1455;
  reg [3-1:0] verilogPut_KeyCollapse_2_1456;
  reg [64-1:0] verilogPut_Data_2_1457;
  reg [64-1:0] verilogPut_Key_3_1458;
  reg [1-1:0] verilogPut_KeyCompares_3_1459;
  reg [3-1:0] verilogPut_KeyCollapse_3_1460;
  reg [64-1:0] verilogPut_Data_3_1461;
  reg [1-1:0] verilogPut_Found_1462;
  reg [64-1:0] verilogPut_Key_1463;
  reg [64-1:0] verilogPut_FoundKey_1464;
  reg [64-1:0] verilogPut_Data_1465;
  reg [4-1:0] verilogPut_BtreeIndex_1466;
  reg [3-1:0] verilogPut_StuckIndex_1467;
  reg [1-1:0] verilogPut_MergeSuccess_1468;
  reg [64-1:0] verilogPut_childKey_1469;
  reg [3-1:0] verilogPut_leftChild_1470;
  reg [3-1:0] verilogPut_rightChild_1471;
  reg [4-1:0] verilogPut_childData_1472;
  reg [4-1:0] verilogPut_indexLeft_1473;
  reg [4-1:0] verilogPut_indexRight_1474;
  reg [64-1:0] verilogPut_midKey_1475;
  reg [1-1:0] verilogPut_success_1476;
  reg [1-1:0] verilogPut_test_1477;
  reg [4-1:0] verilogPut_next_1478;
  reg [4-1:0] verilogPut_root_1479;
  reg [1-1:0] verilogPut_isFree_1480;
  integer verilogPut_pc;
  integer verilogPut_stop;
  integer verilogPut_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      verilogPut_pc <= 0;
      verilogPut_stop <= 0;
      verilogPut_returnCode <= 0;
      verilogPut_index_2 <= 0;
      verilogPut_size_3 <= 0;
      verilogPut_isLeaf_4 <= 0;
      verilogPut_nextFree_5 <= 0;
      verilogPut_Key_0_6 <= 0;
      verilogPut_KeyCompares_0_7 <= 0;
      verilogPut_KeyCollapse_0_8 <= 0;
      verilogPut_Data_0_9 <= 0;
      verilogPut_Key_1_10 <= 0;
      verilogPut_KeyCompares_1_11 <= 0;
      verilogPut_KeyCollapse_1_12 <= 0;
      verilogPut_Data_1_13 <= 0;
      verilogPut_Key_2_14 <= 0;
      verilogPut_KeyCompares_2_15 <= 0;
      verilogPut_KeyCollapse_2_16 <= 0;
      verilogPut_Data_2_17 <= 0;
      verilogPut_Key_3_18 <= 0;
      verilogPut_KeyCompares_3_19 <= 0;
      verilogPut_KeyCollapse_3_20 <= 0;
      verilogPut_Data_3_21 <= 0;
      verilogPut_stuckKeys_1_index_22 <= 0;
      verilogPut_stuckKeys_2_index_23 <= 0;
      verilogPut_stuckKeys_2_value_24 <= 0;
      verilogPut_stuckKeys_2_value_25 <= 0;
      verilogPut_stuckKeys_2_value_26 <= 0;
      verilogPut_stuckKeys_2_value_27 <= 0;
      verilogPut_stuckData_3_index_28 <= 0;
      verilogPut_stuckData_4_index_29 <= 0;
      verilogPut_stuckData_4_value_30 <= 0;
      verilogPut_stuckData_4_value_31 <= 0;
      verilogPut_stuckData_4_value_32 <= 0;
      verilogPut_stuckData_4_value_33 <= 0;
      verilogPut_stuckSize_5_index_34 <= 0;
      verilogPut_stuckSize_6_index_35 <= 0;
      verilogPut_stuckSize_6_value_36 <= 0;
      verilogPut_stuckIsLeaf_7_index_37 <= 0;
      verilogPut_stuckIsLeaf_8_index_38 <= 0;
      verilogPut_stuckIsLeaf_8_value_39 <= 0;
      verilogPut_Found_40 <= 0;
      verilogPut_Key_41 <= 0;
      verilogPut_FoundKey_42 <= 0;
      verilogPut_Data_43 <= 0;
      verilogPut_BtreeIndex_44 <= 0;
      verilogPut_StuckIndex_45 <= 0;
      verilogPut_MergeSuccess_46 <= 0;
      verilogPut_index_47 <= 0;
      verilogPut_size_48 <= 0;
      verilogPut_isLeaf_49 <= 0;
      verilogPut_nextFree_50 <= 0;
      verilogPut_Key_0_51 <= 0;
      verilogPut_KeyCompares_0_52 <= 0;
      verilogPut_KeyCollapse_0_53 <= 0;
      verilogPut_Data_0_54 <= 0;
      verilogPut_Key_1_55 <= 0;
      verilogPut_KeyCompares_1_56 <= 0;
      verilogPut_KeyCollapse_1_57 <= 0;
      verilogPut_Data_1_58 <= 0;
      verilogPut_Key_2_59 <= 0;
      verilogPut_KeyCompares_2_60 <= 0;
      verilogPut_KeyCollapse_2_61 <= 0;
      verilogPut_Data_2_62 <= 0;
      verilogPut_Key_3_63 <= 0;
      verilogPut_KeyCompares_3_64 <= 0;
      verilogPut_KeyCollapse_3_65 <= 0;
      verilogPut_Data_3_66 <= 0;
      verilogPut_Found_67 <= 0;
      verilogPut_Key_68 <= 0;
      verilogPut_FoundKey_69 <= 0;
      verilogPut_Data_70 <= 0;
      verilogPut_BtreeIndex_71 <= 0;
      verilogPut_StuckIndex_72 <= 0;
      verilogPut_MergeSuccess_73 <= 0;
      verilogPut_index_74 <= 0;
      verilogPut_size_75 <= 0;
      verilogPut_isLeaf_76 <= 0;
      verilogPut_nextFree_77 <= 0;
      verilogPut_Key_0_78 <= 0;
      verilogPut_KeyCompares_0_79 <= 0;
      verilogPut_KeyCollapse_0_80 <= 0;
      verilogPut_Data_0_81 <= 0;
      verilogPut_Key_1_82 <= 0;
      verilogPut_KeyCompares_1_83 <= 0;
      verilogPut_KeyCollapse_1_84 <= 0;
      verilogPut_Data_1_85 <= 0;
      verilogPut_Key_2_86 <= 0;
      verilogPut_KeyCompares_2_87 <= 0;
      verilogPut_KeyCollapse_2_88 <= 0;
      verilogPut_Data_2_89 <= 0;
      verilogPut_Key_3_90 <= 0;
      verilogPut_KeyCompares_3_91 <= 0;
      verilogPut_KeyCollapse_3_92 <= 0;
      verilogPut_Data_3_93 <= 0;
      verilogPut_Found_94 <= 0;
      verilogPut_Key_95 <= 0;
      verilogPut_FoundKey_96 <= 0;
      verilogPut_Data_97 <= 0;
      verilogPut_BtreeIndex_98 <= 0;
      verilogPut_StuckIndex_99 <= 0;
      verilogPut_MergeSuccess_100 <= 0;
      verilogPut_child_101 <= 0;
      verilogPut_parent_102 <= 0;
      verilogPut_childInparent_103 <= 0;
      verilogPut_found_104 <= 0;
      verilogPut_full_105 <= 0;
      verilogPut_i_106 <= 0;
      verilogPut_notFull_107 <= 0;
      verilogPut_index_108 <= 0;
      verilogPut_size_109 <= 0;
      verilogPut_isLeaf_110 <= 0;
      verilogPut_nextFree_111 <= 0;
      verilogPut_Key_0_112 <= 0;
      verilogPut_KeyCompares_0_113 <= 0;
      verilogPut_KeyCollapse_0_114 <= 0;
      verilogPut_Data_0_115 <= 0;
      verilogPut_Key_1_116 <= 0;
      verilogPut_KeyCompares_1_117 <= 0;
      verilogPut_KeyCollapse_1_118 <= 0;
      verilogPut_Data_1_119 <= 0;
      verilogPut_Key_2_120 <= 0;
      verilogPut_KeyCompares_2_121 <= 0;
      verilogPut_KeyCollapse_2_122 <= 0;
      verilogPut_Data_2_123 <= 0;
      verilogPut_Key_3_124 <= 0;
      verilogPut_KeyCompares_3_125 <= 0;
      verilogPut_KeyCollapse_3_126 <= 0;
      verilogPut_Data_3_127 <= 0;
      verilogPut_Found_128 <= 0;
      verilogPut_Key_129 <= 0;
      verilogPut_FoundKey_130 <= 0;
      verilogPut_Data_131 <= 0;
      verilogPut_BtreeIndex_132 <= 0;
      verilogPut_StuckIndex_133 <= 0;
      verilogPut_MergeSuccess_134 <= 0;
      verilogPut_index_135 <= 0;
      verilogPut_size_136 <= 0;
      verilogPut_isLeaf_137 <= 0;
      verilogPut_nextFree_138 <= 0;
      verilogPut_Key_0_139 <= 0;
      verilogPut_KeyCompares_0_140 <= 0;
      verilogPut_KeyCollapse_0_141 <= 0;
      verilogPut_Data_0_142 <= 0;
      verilogPut_Key_1_143 <= 0;
      verilogPut_KeyCompares_1_144 <= 0;
      verilogPut_KeyCollapse_1_145 <= 0;
      verilogPut_Data_1_146 <= 0;
      verilogPut_Key_2_147 <= 0;
      verilogPut_KeyCompares_2_148 <= 0;
      verilogPut_KeyCollapse_2_149 <= 0;
      verilogPut_Data_2_150 <= 0;
      verilogPut_Key_3_151 <= 0;
      verilogPut_KeyCompares_3_152 <= 0;
      verilogPut_KeyCollapse_3_153 <= 0;
      verilogPut_Data_3_154 <= 0;
      verilogPut_Found_155 <= 0;
      verilogPut_Key_156 <= 0;
      verilogPut_FoundKey_157 <= 0;
      verilogPut_Data_158 <= 0;
      verilogPut_BtreeIndex_159 <= 0;
      verilogPut_StuckIndex_160 <= 0;
      verilogPut_MergeSuccess_161 <= 0;
      verilogPut_index_162 <= 0;
      verilogPut_size_163 <= 0;
      verilogPut_isLeaf_164 <= 0;
      verilogPut_nextFree_165 <= 0;
      verilogPut_Key_0_166 <= 0;
      verilogPut_KeyCompares_0_167 <= 0;
      verilogPut_KeyCollapse_0_168 <= 0;
      verilogPut_Data_0_169 <= 0;
      verilogPut_Key_1_170 <= 0;
      verilogPut_KeyCompares_1_171 <= 0;
      verilogPut_KeyCollapse_1_172 <= 0;
      verilogPut_Data_1_173 <= 0;
      verilogPut_Key_2_174 <= 0;
      verilogPut_KeyCompares_2_175 <= 0;
      verilogPut_KeyCollapse_2_176 <= 0;
      verilogPut_Data_2_177 <= 0;
      verilogPut_Key_3_178 <= 0;
      verilogPut_KeyCompares_3_179 <= 0;
      verilogPut_KeyCollapse_3_180 <= 0;
      verilogPut_Data_3_181 <= 0;
      verilogPut_Found_182 <= 0;
      verilogPut_Key_183 <= 0;
      verilogPut_FoundKey_184 <= 0;
      verilogPut_Data_185 <= 0;
      verilogPut_BtreeIndex_186 <= 0;
      verilogPut_StuckIndex_187 <= 0;
      verilogPut_MergeSuccess_188 <= 0;
      verilogPut_indexLeft_189 <= 0;
      verilogPut_indexRight_190 <= 0;
      verilogPut_midKey_191 <= 0;
      verilogPut_freeNext_9_index_192 <= 0;
      verilogPut_freeNext_10_index_193 <= 0;
      verilogPut_freeNext_10_value_194 <= 0;
      verilogPut_stuckIsFree_11_index_195 <= 0;
      verilogPut_stuckIsFree_11_value_196 <= 0;
      verilogPut_root_197 <= 0;
      verilogPut_next_198 <= 0;
      verilogPut_isLeaf_199 <= 0;
      verilogPut_isFree_200 <= 0;
      verilogPut_root_201 <= 0;
      verilogPut_next_202 <= 0;
      verilogPut_isLeaf_203 <= 0;
      verilogPut_isFree_204 <= 0;
      verilogPut_i_205 <= 0;
      verilogPut_notFull_206 <= 0;
      verilogPut_index_207 <= 0;
      verilogPut_size_208 <= 0;
      verilogPut_isLeaf_209 <= 0;
      verilogPut_nextFree_210 <= 0;
      verilogPut_Key_0_211 <= 0;
      verilogPut_KeyCompares_0_212 <= 0;
      verilogPut_KeyCollapse_0_213 <= 0;
      verilogPut_Data_0_214 <= 0;
      verilogPut_Key_1_215 <= 0;
      verilogPut_KeyCompares_1_216 <= 0;
      verilogPut_KeyCollapse_1_217 <= 0;
      verilogPut_Data_1_218 <= 0;
      verilogPut_Key_2_219 <= 0;
      verilogPut_KeyCompares_2_220 <= 0;
      verilogPut_KeyCollapse_2_221 <= 0;
      verilogPut_Data_2_222 <= 0;
      verilogPut_Key_3_223 <= 0;
      verilogPut_KeyCompares_3_224 <= 0;
      verilogPut_KeyCollapse_3_225 <= 0;
      verilogPut_Data_3_226 <= 0;
      verilogPut_Found_227 <= 0;
      verilogPut_Key_228 <= 0;
      verilogPut_FoundKey_229 <= 0;
      verilogPut_Data_230 <= 0;
      verilogPut_BtreeIndex_231 <= 0;
      verilogPut_StuckIndex_232 <= 0;
      verilogPut_MergeSuccess_233 <= 0;
      verilogPut_index_234 <= 0;
      verilogPut_size_235 <= 0;
      verilogPut_isLeaf_236 <= 0;
      verilogPut_nextFree_237 <= 0;
      verilogPut_Key_0_238 <= 0;
      verilogPut_KeyCompares_0_239 <= 0;
      verilogPut_KeyCollapse_0_240 <= 0;
      verilogPut_Data_0_241 <= 0;
      verilogPut_Key_1_242 <= 0;
      verilogPut_KeyCompares_1_243 <= 0;
      verilogPut_KeyCollapse_1_244 <= 0;
      verilogPut_Data_1_245 <= 0;
      verilogPut_Key_2_246 <= 0;
      verilogPut_KeyCompares_2_247 <= 0;
      verilogPut_KeyCollapse_2_248 <= 0;
      verilogPut_Data_2_249 <= 0;
      verilogPut_Key_3_250 <= 0;
      verilogPut_KeyCompares_3_251 <= 0;
      verilogPut_KeyCollapse_3_252 <= 0;
      verilogPut_Data_3_253 <= 0;
      verilogPut_Found_254 <= 0;
      verilogPut_Key_255 <= 0;
      verilogPut_FoundKey_256 <= 0;
      verilogPut_Data_257 <= 0;
      verilogPut_BtreeIndex_258 <= 0;
      verilogPut_StuckIndex_259 <= 0;
      verilogPut_MergeSuccess_260 <= 0;
      verilogPut_index_261 <= 0;
      verilogPut_size_262 <= 0;
      verilogPut_isLeaf_263 <= 0;
      verilogPut_nextFree_264 <= 0;
      verilogPut_Key_0_265 <= 0;
      verilogPut_KeyCompares_0_266 <= 0;
      verilogPut_KeyCollapse_0_267 <= 0;
      verilogPut_Data_0_268 <= 0;
      verilogPut_Key_1_269 <= 0;
      verilogPut_KeyCompares_1_270 <= 0;
      verilogPut_KeyCollapse_1_271 <= 0;
      verilogPut_Data_1_272 <= 0;
      verilogPut_Key_2_273 <= 0;
      verilogPut_KeyCompares_2_274 <= 0;
      verilogPut_KeyCollapse_2_275 <= 0;
      verilogPut_Data_2_276 <= 0;
      verilogPut_Key_3_277 <= 0;
      verilogPut_KeyCompares_3_278 <= 0;
      verilogPut_KeyCollapse_3_279 <= 0;
      verilogPut_Data_3_280 <= 0;
      verilogPut_Found_281 <= 0;
      verilogPut_Key_282 <= 0;
      verilogPut_FoundKey_283 <= 0;
      verilogPut_Data_284 <= 0;
      verilogPut_BtreeIndex_285 <= 0;
      verilogPut_StuckIndex_286 <= 0;
      verilogPut_MergeSuccess_287 <= 0;
      verilogPut_indexLeft_288 <= 0;
      verilogPut_indexRight_289 <= 0;
      verilogPut_midKey_290 <= 0;
      verilogPut_root_291 <= 0;
      verilogPut_next_292 <= 0;
      verilogPut_isLeaf_293 <= 0;
      verilogPut_isFree_294 <= 0;
      verilogPut_root_295 <= 0;
      verilogPut_next_296 <= 0;
      verilogPut_isLeaf_297 <= 0;
      verilogPut_isFree_298 <= 0;
      verilogPut_index_299 <= 0;
      verilogPut_size_300 <= 0;
      verilogPut_isLeaf_301 <= 0;
      verilogPut_nextFree_302 <= 0;
      verilogPut_Key_0_303 <= 0;
      verilogPut_KeyCompares_0_304 <= 0;
      verilogPut_KeyCollapse_0_305 <= 0;
      verilogPut_Data_0_306 <= 0;
      verilogPut_Key_1_307 <= 0;
      verilogPut_KeyCompares_1_308 <= 0;
      verilogPut_KeyCollapse_1_309 <= 0;
      verilogPut_Data_1_310 <= 0;
      verilogPut_Key_2_311 <= 0;
      verilogPut_KeyCompares_2_312 <= 0;
      verilogPut_KeyCollapse_2_313 <= 0;
      verilogPut_Data_2_314 <= 0;
      verilogPut_Key_3_315 <= 0;
      verilogPut_KeyCompares_3_316 <= 0;
      verilogPut_KeyCollapse_3_317 <= 0;
      verilogPut_Data_3_318 <= 0;
      verilogPut_Found_319 <= 0;
      verilogPut_Key_320 <= 0;
      verilogPut_FoundKey_321 <= 0;
      verilogPut_Data_322 <= 0;
      verilogPut_BtreeIndex_323 <= 0;
      verilogPut_StuckIndex_324 <= 0;
      verilogPut_MergeSuccess_325 <= 0;
      verilogPut_index_326 <= 0;
      verilogPut_size_327 <= 0;
      verilogPut_isLeaf_328 <= 0;
      verilogPut_nextFree_329 <= 0;
      verilogPut_Key_0_330 <= 0;
      verilogPut_KeyCompares_0_331 <= 0;
      verilogPut_KeyCollapse_0_332 <= 0;
      verilogPut_Data_0_333 <= 0;
      verilogPut_Key_1_334 <= 0;
      verilogPut_KeyCompares_1_335 <= 0;
      verilogPut_KeyCollapse_1_336 <= 0;
      verilogPut_Data_1_337 <= 0;
      verilogPut_Key_2_338 <= 0;
      verilogPut_KeyCompares_2_339 <= 0;
      verilogPut_KeyCollapse_2_340 <= 0;
      verilogPut_Data_2_341 <= 0;
      verilogPut_Key_3_342 <= 0;
      verilogPut_KeyCompares_3_343 <= 0;
      verilogPut_KeyCollapse_3_344 <= 0;
      verilogPut_Data_3_345 <= 0;
      verilogPut_Found_346 <= 0;
      verilogPut_Key_347 <= 0;
      verilogPut_FoundKey_348 <= 0;
      verilogPut_Data_349 <= 0;
      verilogPut_BtreeIndex_350 <= 0;
      verilogPut_StuckIndex_351 <= 0;
      verilogPut_MergeSuccess_352 <= 0;
      verilogPut_index_353 <= 0;
      verilogPut_size_354 <= 0;
      verilogPut_isLeaf_355 <= 0;
      verilogPut_nextFree_356 <= 0;
      verilogPut_Key_0_357 <= 0;
      verilogPut_KeyCompares_0_358 <= 0;
      verilogPut_KeyCollapse_0_359 <= 0;
      verilogPut_Data_0_360 <= 0;
      verilogPut_Key_1_361 <= 0;
      verilogPut_KeyCompares_1_362 <= 0;
      verilogPut_KeyCollapse_1_363 <= 0;
      verilogPut_Data_1_364 <= 0;
      verilogPut_Key_2_365 <= 0;
      verilogPut_KeyCompares_2_366 <= 0;
      verilogPut_KeyCollapse_2_367 <= 0;
      verilogPut_Data_2_368 <= 0;
      verilogPut_Key_3_369 <= 0;
      verilogPut_KeyCompares_3_370 <= 0;
      verilogPut_KeyCollapse_3_371 <= 0;
      verilogPut_Data_3_372 <= 0;
      verilogPut_Found_373 <= 0;
      verilogPut_Key_374 <= 0;
      verilogPut_FoundKey_375 <= 0;
      verilogPut_Data_376 <= 0;
      verilogPut_BtreeIndex_377 <= 0;
      verilogPut_StuckIndex_378 <= 0;
      verilogPut_MergeSuccess_379 <= 0;
      verilogPut_index_380 <= 0;
      verilogPut_size_381 <= 0;
      verilogPut_isLeaf_382 <= 0;
      verilogPut_nextFree_383 <= 0;
      verilogPut_Key_0_384 <= 0;
      verilogPut_KeyCompares_0_385 <= 0;
      verilogPut_KeyCollapse_0_386 <= 0;
      verilogPut_Data_0_387 <= 0;
      verilogPut_Key_1_388 <= 0;
      verilogPut_KeyCompares_1_389 <= 0;
      verilogPut_KeyCollapse_1_390 <= 0;
      verilogPut_Data_1_391 <= 0;
      verilogPut_Key_2_392 <= 0;
      verilogPut_KeyCompares_2_393 <= 0;
      verilogPut_KeyCollapse_2_394 <= 0;
      verilogPut_Data_2_395 <= 0;
      verilogPut_Key_3_396 <= 0;
      verilogPut_KeyCompares_3_397 <= 0;
      verilogPut_KeyCollapse_3_398 <= 0;
      verilogPut_Data_3_399 <= 0;
      verilogPut_Found_400 <= 0;
      verilogPut_Key_401 <= 0;
      verilogPut_FoundKey_402 <= 0;
      verilogPut_Data_403 <= 0;
      verilogPut_BtreeIndex_404 <= 0;
      verilogPut_StuckIndex_405 <= 0;
      verilogPut_MergeSuccess_406 <= 0;
      verilogPut_childKey_407 <= 0;
      verilogPut_childData_408 <= 0;
      verilogPut_indexLeft_409 <= 0;
      verilogPut_indexRight_410 <= 0;
      verilogPut_midKey_411 <= 0;
      verilogPut_root_412 <= 0;
      verilogPut_next_413 <= 0;
      verilogPut_isLeaf_414 <= 0;
      verilogPut_isFree_415 <= 0;
      verilogPut_index_416 <= 0;
      verilogPut_size_417 <= 0;
      verilogPut_isLeaf_418 <= 0;
      verilogPut_nextFree_419 <= 0;
      verilogPut_Key_0_420 <= 0;
      verilogPut_KeyCompares_0_421 <= 0;
      verilogPut_KeyCollapse_0_422 <= 0;
      verilogPut_Data_0_423 <= 0;
      verilogPut_Key_1_424 <= 0;
      verilogPut_KeyCompares_1_425 <= 0;
      verilogPut_KeyCollapse_1_426 <= 0;
      verilogPut_Data_1_427 <= 0;
      verilogPut_Key_2_428 <= 0;
      verilogPut_KeyCompares_2_429 <= 0;
      verilogPut_KeyCollapse_2_430 <= 0;
      verilogPut_Data_2_431 <= 0;
      verilogPut_Key_3_432 <= 0;
      verilogPut_KeyCompares_3_433 <= 0;
      verilogPut_KeyCollapse_3_434 <= 0;
      verilogPut_Data_3_435 <= 0;
      verilogPut_Found_436 <= 0;
      verilogPut_Key_437 <= 0;
      verilogPut_FoundKey_438 <= 0;
      verilogPut_Data_439 <= 0;
      verilogPut_BtreeIndex_440 <= 0;
      verilogPut_StuckIndex_441 <= 0;
      verilogPut_MergeSuccess_442 <= 0;
      verilogPut_index_443 <= 0;
      verilogPut_size_444 <= 0;
      verilogPut_isLeaf_445 <= 0;
      verilogPut_nextFree_446 <= 0;
      verilogPut_Key_0_447 <= 0;
      verilogPut_KeyCompares_0_448 <= 0;
      verilogPut_KeyCollapse_0_449 <= 0;
      verilogPut_Data_0_450 <= 0;
      verilogPut_Key_1_451 <= 0;
      verilogPut_KeyCompares_1_452 <= 0;
      verilogPut_KeyCollapse_1_453 <= 0;
      verilogPut_Data_1_454 <= 0;
      verilogPut_Key_2_455 <= 0;
      verilogPut_KeyCompares_2_456 <= 0;
      verilogPut_KeyCollapse_2_457 <= 0;
      verilogPut_Data_2_458 <= 0;
      verilogPut_Key_3_459 <= 0;
      verilogPut_KeyCompares_3_460 <= 0;
      verilogPut_KeyCollapse_3_461 <= 0;
      verilogPut_Data_3_462 <= 0;
      verilogPut_Found_463 <= 0;
      verilogPut_Key_464 <= 0;
      verilogPut_FoundKey_465 <= 0;
      verilogPut_Data_466 <= 0;
      verilogPut_BtreeIndex_467 <= 0;
      verilogPut_StuckIndex_468 <= 0;
      verilogPut_MergeSuccess_469 <= 0;
      verilogPut_index_470 <= 0;
      verilogPut_size_471 <= 0;
      verilogPut_isLeaf_472 <= 0;
      verilogPut_nextFree_473 <= 0;
      verilogPut_Key_0_474 <= 0;
      verilogPut_KeyCompares_0_475 <= 0;
      verilogPut_KeyCollapse_0_476 <= 0;
      verilogPut_Data_0_477 <= 0;
      verilogPut_Key_1_478 <= 0;
      verilogPut_KeyCompares_1_479 <= 0;
      verilogPut_KeyCollapse_1_480 <= 0;
      verilogPut_Data_1_481 <= 0;
      verilogPut_Key_2_482 <= 0;
      verilogPut_KeyCompares_2_483 <= 0;
      verilogPut_KeyCollapse_2_484 <= 0;
      verilogPut_Data_2_485 <= 0;
      verilogPut_Key_3_486 <= 0;
      verilogPut_KeyCompares_3_487 <= 0;
      verilogPut_KeyCollapse_3_488 <= 0;
      verilogPut_Data_3_489 <= 0;
      verilogPut_Found_490 <= 0;
      verilogPut_Key_491 <= 0;
      verilogPut_FoundKey_492 <= 0;
      verilogPut_Data_493 <= 0;
      verilogPut_BtreeIndex_494 <= 0;
      verilogPut_StuckIndex_495 <= 0;
      verilogPut_MergeSuccess_496 <= 0;
      verilogPut_childIndex_497 <= 0;
      verilogPut_leftIndex_498 <= 0;
      verilogPut_midKey_499 <= 0;
      verilogPut_root_500 <= 0;
      verilogPut_next_501 <= 0;
      verilogPut_isLeaf_502 <= 0;
      verilogPut_isFree_503 <= 0;
      verilogPut_i_504 <= 0;
      verilogPut_notFull_505 <= 0;
      verilogPut_index_506 <= 0;
      verilogPut_size_507 <= 0;
      verilogPut_isLeaf_508 <= 0;
      verilogPut_nextFree_509 <= 0;
      verilogPut_Key_0_510 <= 0;
      verilogPut_KeyCompares_0_511 <= 0;
      verilogPut_KeyCollapse_0_512 <= 0;
      verilogPut_Data_0_513 <= 0;
      verilogPut_Key_1_514 <= 0;
      verilogPut_KeyCompares_1_515 <= 0;
      verilogPut_KeyCollapse_1_516 <= 0;
      verilogPut_Data_1_517 <= 0;
      verilogPut_Key_2_518 <= 0;
      verilogPut_KeyCompares_2_519 <= 0;
      verilogPut_KeyCollapse_2_520 <= 0;
      verilogPut_Data_2_521 <= 0;
      verilogPut_Key_3_522 <= 0;
      verilogPut_KeyCompares_3_523 <= 0;
      verilogPut_KeyCollapse_3_524 <= 0;
      verilogPut_Data_3_525 <= 0;
      verilogPut_Found_526 <= 0;
      verilogPut_Key_527 <= 0;
      verilogPut_FoundKey_528 <= 0;
      verilogPut_Data_529 <= 0;
      verilogPut_BtreeIndex_530 <= 0;
      verilogPut_StuckIndex_531 <= 0;
      verilogPut_MergeSuccess_532 <= 0;
      verilogPut_index_533 <= 0;
      verilogPut_size_534 <= 0;
      verilogPut_isLeaf_535 <= 0;
      verilogPut_nextFree_536 <= 0;
      verilogPut_Key_0_537 <= 0;
      verilogPut_KeyCompares_0_538 <= 0;
      verilogPut_KeyCollapse_0_539 <= 0;
      verilogPut_Data_0_540 <= 0;
      verilogPut_Key_1_541 <= 0;
      verilogPut_KeyCompares_1_542 <= 0;
      verilogPut_KeyCollapse_1_543 <= 0;
      verilogPut_Data_1_544 <= 0;
      verilogPut_Key_2_545 <= 0;
      verilogPut_KeyCompares_2_546 <= 0;
      verilogPut_KeyCollapse_2_547 <= 0;
      verilogPut_Data_2_548 <= 0;
      verilogPut_Key_3_549 <= 0;
      verilogPut_KeyCompares_3_550 <= 0;
      verilogPut_KeyCollapse_3_551 <= 0;
      verilogPut_Data_3_552 <= 0;
      verilogPut_Found_553 <= 0;
      verilogPut_Key_554 <= 0;
      verilogPut_FoundKey_555 <= 0;
      verilogPut_Data_556 <= 0;
      verilogPut_BtreeIndex_557 <= 0;
      verilogPut_StuckIndex_558 <= 0;
      verilogPut_MergeSuccess_559 <= 0;
      verilogPut_index_560 <= 0;
      verilogPut_size_561 <= 0;
      verilogPut_isLeaf_562 <= 0;
      verilogPut_nextFree_563 <= 0;
      verilogPut_Key_0_564 <= 0;
      verilogPut_KeyCompares_0_565 <= 0;
      verilogPut_KeyCollapse_0_566 <= 0;
      verilogPut_Data_0_567 <= 0;
      verilogPut_Key_1_568 <= 0;
      verilogPut_KeyCompares_1_569 <= 0;
      verilogPut_KeyCollapse_1_570 <= 0;
      verilogPut_Data_1_571 <= 0;
      verilogPut_Key_2_572 <= 0;
      verilogPut_KeyCompares_2_573 <= 0;
      verilogPut_KeyCollapse_2_574 <= 0;
      verilogPut_Data_2_575 <= 0;
      verilogPut_Key_3_576 <= 0;
      verilogPut_KeyCompares_3_577 <= 0;
      verilogPut_KeyCollapse_3_578 <= 0;
      verilogPut_Data_3_579 <= 0;
      verilogPut_Found_580 <= 0;
      verilogPut_Key_581 <= 0;
      verilogPut_FoundKey_582 <= 0;
      verilogPut_Data_583 <= 0;
      verilogPut_BtreeIndex_584 <= 0;
      verilogPut_StuckIndex_585 <= 0;
      verilogPut_MergeSuccess_586 <= 0;
      verilogPut_index_587 <= 0;
      verilogPut_size_588 <= 0;
      verilogPut_isLeaf_589 <= 0;
      verilogPut_nextFree_590 <= 0;
      verilogPut_Key_0_591 <= 0;
      verilogPut_KeyCompares_0_592 <= 0;
      verilogPut_KeyCollapse_0_593 <= 0;
      verilogPut_Data_0_594 <= 0;
      verilogPut_Key_1_595 <= 0;
      verilogPut_KeyCompares_1_596 <= 0;
      verilogPut_KeyCollapse_1_597 <= 0;
      verilogPut_Data_1_598 <= 0;
      verilogPut_Key_2_599 <= 0;
      verilogPut_KeyCompares_2_600 <= 0;
      verilogPut_KeyCollapse_2_601 <= 0;
      verilogPut_Data_2_602 <= 0;
      verilogPut_Key_3_603 <= 0;
      verilogPut_KeyCompares_3_604 <= 0;
      verilogPut_KeyCollapse_3_605 <= 0;
      verilogPut_Data_3_606 <= 0;
      verilogPut_Found_607 <= 0;
      verilogPut_Key_608 <= 0;
      verilogPut_FoundKey_609 <= 0;
      verilogPut_Data_610 <= 0;
      verilogPut_BtreeIndex_611 <= 0;
      verilogPut_StuckIndex_612 <= 0;
      verilogPut_MergeSuccess_613 <= 0;
      verilogPut_childKey_614 <= 0;
      verilogPut_childData_615 <= 0;
      verilogPut_indexLeft_616 <= 0;
      verilogPut_indexRight_617 <= 0;
      verilogPut_midKey_618 <= 0;
      verilogPut_root_619 <= 0;
      verilogPut_next_620 <= 0;
      verilogPut_isLeaf_621 <= 0;
      verilogPut_isFree_622 <= 0;
      verilogPut_index_623 <= 0;
      verilogPut_size_624 <= 0;
      verilogPut_isLeaf_625 <= 0;
      verilogPut_nextFree_626 <= 0;
      verilogPut_Key_0_627 <= 0;
      verilogPut_KeyCompares_0_628 <= 0;
      verilogPut_KeyCollapse_0_629 <= 0;
      verilogPut_Data_0_630 <= 0;
      verilogPut_Key_1_631 <= 0;
      verilogPut_KeyCompares_1_632 <= 0;
      verilogPut_KeyCollapse_1_633 <= 0;
      verilogPut_Data_1_634 <= 0;
      verilogPut_Key_2_635 <= 0;
      verilogPut_KeyCompares_2_636 <= 0;
      verilogPut_KeyCollapse_2_637 <= 0;
      verilogPut_Data_2_638 <= 0;
      verilogPut_Key_3_639 <= 0;
      verilogPut_KeyCompares_3_640 <= 0;
      verilogPut_KeyCollapse_3_641 <= 0;
      verilogPut_Data_3_642 <= 0;
      verilogPut_Found_643 <= 0;
      verilogPut_Key_644 <= 0;
      verilogPut_FoundKey_645 <= 0;
      verilogPut_Data_646 <= 0;
      verilogPut_BtreeIndex_647 <= 0;
      verilogPut_StuckIndex_648 <= 0;
      verilogPut_MergeSuccess_649 <= 0;
      verilogPut_index_650 <= 0;
      verilogPut_size_651 <= 0;
      verilogPut_isLeaf_652 <= 0;
      verilogPut_nextFree_653 <= 0;
      verilogPut_Key_0_654 <= 0;
      verilogPut_KeyCompares_0_655 <= 0;
      verilogPut_KeyCollapse_0_656 <= 0;
      verilogPut_Data_0_657 <= 0;
      verilogPut_Key_1_658 <= 0;
      verilogPut_KeyCompares_1_659 <= 0;
      verilogPut_KeyCollapse_1_660 <= 0;
      verilogPut_Data_1_661 <= 0;
      verilogPut_Key_2_662 <= 0;
      verilogPut_KeyCompares_2_663 <= 0;
      verilogPut_KeyCollapse_2_664 <= 0;
      verilogPut_Data_2_665 <= 0;
      verilogPut_Key_3_666 <= 0;
      verilogPut_KeyCompares_3_667 <= 0;
      verilogPut_KeyCollapse_3_668 <= 0;
      verilogPut_Data_3_669 <= 0;
      verilogPut_Found_670 <= 0;
      verilogPut_Key_671 <= 0;
      verilogPut_FoundKey_672 <= 0;
      verilogPut_Data_673 <= 0;
      verilogPut_BtreeIndex_674 <= 0;
      verilogPut_StuckIndex_675 <= 0;
      verilogPut_MergeSuccess_676 <= 0;
      verilogPut_index_677 <= 0;
      verilogPut_size_678 <= 0;
      verilogPut_isLeaf_679 <= 0;
      verilogPut_nextFree_680 <= 0;
      verilogPut_Key_0_681 <= 0;
      verilogPut_KeyCompares_0_682 <= 0;
      verilogPut_KeyCollapse_0_683 <= 0;
      verilogPut_Data_0_684 <= 0;
      verilogPut_Key_1_685 <= 0;
      verilogPut_KeyCompares_1_686 <= 0;
      verilogPut_KeyCollapse_1_687 <= 0;
      verilogPut_Data_1_688 <= 0;
      verilogPut_Key_2_689 <= 0;
      verilogPut_KeyCompares_2_690 <= 0;
      verilogPut_KeyCollapse_2_691 <= 0;
      verilogPut_Data_2_692 <= 0;
      verilogPut_Key_3_693 <= 0;
      verilogPut_KeyCompares_3_694 <= 0;
      verilogPut_KeyCollapse_3_695 <= 0;
      verilogPut_Data_3_696 <= 0;
      verilogPut_Found_697 <= 0;
      verilogPut_Key_698 <= 0;
      verilogPut_FoundKey_699 <= 0;
      verilogPut_Data_700 <= 0;
      verilogPut_BtreeIndex_701 <= 0;
      verilogPut_StuckIndex_702 <= 0;
      verilogPut_MergeSuccess_703 <= 0;
      verilogPut_index_704 <= 0;
      verilogPut_size_705 <= 0;
      verilogPut_isLeaf_706 <= 0;
      verilogPut_nextFree_707 <= 0;
      verilogPut_Key_0_708 <= 0;
      verilogPut_KeyCompares_0_709 <= 0;
      verilogPut_KeyCollapse_0_710 <= 0;
      verilogPut_Data_0_711 <= 0;
      verilogPut_Key_1_712 <= 0;
      verilogPut_KeyCompares_1_713 <= 0;
      verilogPut_KeyCollapse_1_714 <= 0;
      verilogPut_Data_1_715 <= 0;
      verilogPut_Key_2_716 <= 0;
      verilogPut_KeyCompares_2_717 <= 0;
      verilogPut_KeyCollapse_2_718 <= 0;
      verilogPut_Data_2_719 <= 0;
      verilogPut_Key_3_720 <= 0;
      verilogPut_KeyCompares_3_721 <= 0;
      verilogPut_KeyCollapse_3_722 <= 0;
      verilogPut_Data_3_723 <= 0;
      verilogPut_Found_724 <= 0;
      verilogPut_Key_725 <= 0;
      verilogPut_FoundKey_726 <= 0;
      verilogPut_Data_727 <= 0;
      verilogPut_BtreeIndex_728 <= 0;
      verilogPut_StuckIndex_729 <= 0;
      verilogPut_MergeSuccess_730 <= 0;
      verilogPut_childKey_731 <= 0;
      verilogPut_childData_732 <= 0;
      verilogPut_indexLeft_733 <= 0;
      verilogPut_indexRight_734 <= 0;
      verilogPut_midKey_735 <= 0;
      verilogPut_root_736 <= 0;
      verilogPut_next_737 <= 0;
      verilogPut_isLeaf_738 <= 0;
      verilogPut_isFree_739 <= 0;
      verilogPut_index_740 <= 0;
      verilogPut_size_741 <= 0;
      verilogPut_isLeaf_742 <= 0;
      verilogPut_nextFree_743 <= 0;
      verilogPut_Key_0_744 <= 0;
      verilogPut_KeyCompares_0_745 <= 0;
      verilogPut_KeyCollapse_0_746 <= 0;
      verilogPut_Data_0_747 <= 0;
      verilogPut_Key_1_748 <= 0;
      verilogPut_KeyCompares_1_749 <= 0;
      verilogPut_KeyCollapse_1_750 <= 0;
      verilogPut_Data_1_751 <= 0;
      verilogPut_Key_2_752 <= 0;
      verilogPut_KeyCompares_2_753 <= 0;
      verilogPut_KeyCollapse_2_754 <= 0;
      verilogPut_Data_2_755 <= 0;
      verilogPut_Key_3_756 <= 0;
      verilogPut_KeyCompares_3_757 <= 0;
      verilogPut_KeyCollapse_3_758 <= 0;
      verilogPut_Data_3_759 <= 0;
      verilogPut_Found_760 <= 0;
      verilogPut_Key_761 <= 0;
      verilogPut_FoundKey_762 <= 0;
      verilogPut_Data_763 <= 0;
      verilogPut_BtreeIndex_764 <= 0;
      verilogPut_StuckIndex_765 <= 0;
      verilogPut_MergeSuccess_766 <= 0;
      verilogPut_position_767 <= 0;
      verilogPut_index_768 <= 0;
      verilogPut_within_769 <= 0;
      verilogPut_isLeaf_770 <= 0;
      verilogPut_index_771 <= 0;
      verilogPut_size_772 <= 0;
      verilogPut_isLeaf_773 <= 0;
      verilogPut_nextFree_774 <= 0;
      verilogPut_Key_0_775 <= 0;
      verilogPut_KeyCompares_0_776 <= 0;
      verilogPut_KeyCollapse_0_777 <= 0;
      verilogPut_Data_0_778 <= 0;
      verilogPut_Key_1_779 <= 0;
      verilogPut_KeyCompares_1_780 <= 0;
      verilogPut_KeyCollapse_1_781 <= 0;
      verilogPut_Data_1_782 <= 0;
      verilogPut_Key_2_783 <= 0;
      verilogPut_KeyCompares_2_784 <= 0;
      verilogPut_KeyCollapse_2_785 <= 0;
      verilogPut_Data_2_786 <= 0;
      verilogPut_Key_3_787 <= 0;
      verilogPut_KeyCompares_3_788 <= 0;
      verilogPut_KeyCollapse_3_789 <= 0;
      verilogPut_Data_3_790 <= 0;
      verilogPut_Found_791 <= 0;
      verilogPut_Key_792 <= 0;
      verilogPut_FoundKey_793 <= 0;
      verilogPut_Data_794 <= 0;
      verilogPut_BtreeIndex_795 <= 0;
      verilogPut_StuckIndex_796 <= 0;
      verilogPut_MergeSuccess_797 <= 0;
      verilogPut_index_798 <= 0;
      verilogPut_size_799 <= 0;
      verilogPut_isLeaf_800 <= 0;
      verilogPut_nextFree_801 <= 0;
      verilogPut_Key_0_802 <= 0;
      verilogPut_KeyCompares_0_803 <= 0;
      verilogPut_KeyCollapse_0_804 <= 0;
      verilogPut_Data_0_805 <= 0;
      verilogPut_Key_1_806 <= 0;
      verilogPut_KeyCompares_1_807 <= 0;
      verilogPut_KeyCollapse_1_808 <= 0;
      verilogPut_Data_1_809 <= 0;
      verilogPut_Key_2_810 <= 0;
      verilogPut_KeyCompares_2_811 <= 0;
      verilogPut_KeyCollapse_2_812 <= 0;
      verilogPut_Data_2_813 <= 0;
      verilogPut_Key_3_814 <= 0;
      verilogPut_KeyCompares_3_815 <= 0;
      verilogPut_KeyCollapse_3_816 <= 0;
      verilogPut_Data_3_817 <= 0;
      verilogPut_Found_818 <= 0;
      verilogPut_Key_819 <= 0;
      verilogPut_FoundKey_820 <= 0;
      verilogPut_Data_821 <= 0;
      verilogPut_BtreeIndex_822 <= 0;
      verilogPut_StuckIndex_823 <= 0;
      verilogPut_MergeSuccess_824 <= 0;
      verilogPut_index_825 <= 0;
      verilogPut_size_826 <= 0;
      verilogPut_isLeaf_827 <= 0;
      verilogPut_nextFree_828 <= 0;
      verilogPut_Key_0_829 <= 0;
      verilogPut_KeyCompares_0_830 <= 0;
      verilogPut_KeyCollapse_0_831 <= 0;
      verilogPut_Data_0_832 <= 0;
      verilogPut_Key_1_833 <= 0;
      verilogPut_KeyCompares_1_834 <= 0;
      verilogPut_KeyCollapse_1_835 <= 0;
      verilogPut_Data_1_836 <= 0;
      verilogPut_Key_2_837 <= 0;
      verilogPut_KeyCompares_2_838 <= 0;
      verilogPut_KeyCollapse_2_839 <= 0;
      verilogPut_Data_2_840 <= 0;
      verilogPut_Key_3_841 <= 0;
      verilogPut_KeyCompares_3_842 <= 0;
      verilogPut_KeyCollapse_3_843 <= 0;
      verilogPut_Data_3_844 <= 0;
      verilogPut_Found_845 <= 0;
      verilogPut_Key_846 <= 0;
      verilogPut_FoundKey_847 <= 0;
      verilogPut_Data_848 <= 0;
      verilogPut_BtreeIndex_849 <= 0;
      verilogPut_StuckIndex_850 <= 0;
      verilogPut_MergeSuccess_851 <= 0;
      verilogPut_childKey_852 <= 0;
      verilogPut_childData_853 <= 0;
      verilogPut_indexLeft_854 <= 0;
      verilogPut_indexRight_855 <= 0;
      verilogPut_midKey_856 <= 0;
      verilogPut_success_857 <= 0;
      verilogPut_test_858 <= 0;
      verilogPut_next_859 <= 0;
      verilogPut_root_860 <= 0;
      verilogPut_isFree_861 <= 0;
      verilogPut_next_862 <= 0;
      verilogPut_root_863 <= 0;
      verilogPut_isFree_864 <= 0;
      verilogPut_index_865 <= 0;
      verilogPut_size_866 <= 0;
      verilogPut_isLeaf_867 <= 0;
      verilogPut_nextFree_868 <= 0;
      verilogPut_Key_0_869 <= 0;
      verilogPut_KeyCompares_0_870 <= 0;
      verilogPut_KeyCollapse_0_871 <= 0;
      verilogPut_Data_0_872 <= 0;
      verilogPut_Key_1_873 <= 0;
      verilogPut_KeyCompares_1_874 <= 0;
      verilogPut_KeyCollapse_1_875 <= 0;
      verilogPut_Data_1_876 <= 0;
      verilogPut_Key_2_877 <= 0;
      verilogPut_KeyCompares_2_878 <= 0;
      verilogPut_KeyCollapse_2_879 <= 0;
      verilogPut_Data_2_880 <= 0;
      verilogPut_Key_3_881 <= 0;
      verilogPut_KeyCompares_3_882 <= 0;
      verilogPut_KeyCollapse_3_883 <= 0;
      verilogPut_Data_3_884 <= 0;
      verilogPut_Found_885 <= 0;
      verilogPut_Key_886 <= 0;
      verilogPut_FoundKey_887 <= 0;
      verilogPut_Data_888 <= 0;
      verilogPut_BtreeIndex_889 <= 0;
      verilogPut_StuckIndex_890 <= 0;
      verilogPut_MergeSuccess_891 <= 0;
      verilogPut_index_892 <= 0;
      verilogPut_size_893 <= 0;
      verilogPut_isLeaf_894 <= 0;
      verilogPut_nextFree_895 <= 0;
      verilogPut_Key_0_896 <= 0;
      verilogPut_KeyCompares_0_897 <= 0;
      verilogPut_KeyCollapse_0_898 <= 0;
      verilogPut_Data_0_899 <= 0;
      verilogPut_Key_1_900 <= 0;
      verilogPut_KeyCompares_1_901 <= 0;
      verilogPut_KeyCollapse_1_902 <= 0;
      verilogPut_Data_1_903 <= 0;
      verilogPut_Key_2_904 <= 0;
      verilogPut_KeyCompares_2_905 <= 0;
      verilogPut_KeyCollapse_2_906 <= 0;
      verilogPut_Data_2_907 <= 0;
      verilogPut_Key_3_908 <= 0;
      verilogPut_KeyCompares_3_909 <= 0;
      verilogPut_KeyCollapse_3_910 <= 0;
      verilogPut_Data_3_911 <= 0;
      verilogPut_Found_912 <= 0;
      verilogPut_Key_913 <= 0;
      verilogPut_FoundKey_914 <= 0;
      verilogPut_Data_915 <= 0;
      verilogPut_BtreeIndex_916 <= 0;
      verilogPut_StuckIndex_917 <= 0;
      verilogPut_MergeSuccess_918 <= 0;
      verilogPut_index_919 <= 0;
      verilogPut_size_920 <= 0;
      verilogPut_isLeaf_921 <= 0;
      verilogPut_nextFree_922 <= 0;
      verilogPut_Key_0_923 <= 0;
      verilogPut_KeyCompares_0_924 <= 0;
      verilogPut_KeyCollapse_0_925 <= 0;
      verilogPut_Data_0_926 <= 0;
      verilogPut_Key_1_927 <= 0;
      verilogPut_KeyCompares_1_928 <= 0;
      verilogPut_KeyCollapse_1_929 <= 0;
      verilogPut_Data_1_930 <= 0;
      verilogPut_Key_2_931 <= 0;
      verilogPut_KeyCompares_2_932 <= 0;
      verilogPut_KeyCollapse_2_933 <= 0;
      verilogPut_Data_2_934 <= 0;
      verilogPut_Key_3_935 <= 0;
      verilogPut_KeyCompares_3_936 <= 0;
      verilogPut_KeyCollapse_3_937 <= 0;
      verilogPut_Data_3_938 <= 0;
      verilogPut_Found_939 <= 0;
      verilogPut_Key_940 <= 0;
      verilogPut_FoundKey_941 <= 0;
      verilogPut_Data_942 <= 0;
      verilogPut_BtreeIndex_943 <= 0;
      verilogPut_StuckIndex_944 <= 0;
      verilogPut_MergeSuccess_945 <= 0;
      verilogPut_childKey_946 <= 0;
      verilogPut_leftChild_947 <= 0;
      verilogPut_rightChild_948 <= 0;
      verilogPut_childData_949 <= 0;
      verilogPut_indexLeft_950 <= 0;
      verilogPut_indexRight_951 <= 0;
      verilogPut_midKey_952 <= 0;
      verilogPut_success_953 <= 0;
      verilogPut_test_954 <= 0;
      verilogPut_next_955 <= 0;
      verilogPut_root_956 <= 0;
      verilogPut_isFree_957 <= 0;
      verilogPut_next_958 <= 0;
      verilogPut_root_959 <= 0;
      verilogPut_isFree_960 <= 0;
      verilogPut_index_961 <= 0;
      verilogPut_size_962 <= 0;
      verilogPut_isLeaf_963 <= 0;
      verilogPut_nextFree_964 <= 0;
      verilogPut_Key_0_965 <= 0;
      verilogPut_KeyCompares_0_966 <= 0;
      verilogPut_KeyCollapse_0_967 <= 0;
      verilogPut_Data_0_968 <= 0;
      verilogPut_Key_1_969 <= 0;
      verilogPut_KeyCompares_1_970 <= 0;
      verilogPut_KeyCollapse_1_971 <= 0;
      verilogPut_Data_1_972 <= 0;
      verilogPut_Key_2_973 <= 0;
      verilogPut_KeyCompares_2_974 <= 0;
      verilogPut_KeyCollapse_2_975 <= 0;
      verilogPut_Data_2_976 <= 0;
      verilogPut_Key_3_977 <= 0;
      verilogPut_KeyCompares_3_978 <= 0;
      verilogPut_KeyCollapse_3_979 <= 0;
      verilogPut_Data_3_980 <= 0;
      verilogPut_Found_981 <= 0;
      verilogPut_Key_982 <= 0;
      verilogPut_FoundKey_983 <= 0;
      verilogPut_Data_984 <= 0;
      verilogPut_BtreeIndex_985 <= 0;
      verilogPut_StuckIndex_986 <= 0;
      verilogPut_MergeSuccess_987 <= 0;
      verilogPut_index_988 <= 0;
      verilogPut_size_989 <= 0;
      verilogPut_isLeaf_990 <= 0;
      verilogPut_nextFree_991 <= 0;
      verilogPut_Key_0_992 <= 0;
      verilogPut_KeyCompares_0_993 <= 0;
      verilogPut_KeyCollapse_0_994 <= 0;
      verilogPut_Data_0_995 <= 0;
      verilogPut_Key_1_996 <= 0;
      verilogPut_KeyCompares_1_997 <= 0;
      verilogPut_KeyCollapse_1_998 <= 0;
      verilogPut_Data_1_999 <= 0;
      verilogPut_Key_2_1000 <= 0;
      verilogPut_KeyCompares_2_1001 <= 0;
      verilogPut_KeyCollapse_2_1002 <= 0;
      verilogPut_Data_2_1003 <= 0;
      verilogPut_Key_3_1004 <= 0;
      verilogPut_KeyCompares_3_1005 <= 0;
      verilogPut_KeyCollapse_3_1006 <= 0;
      verilogPut_Data_3_1007 <= 0;
      verilogPut_Found_1008 <= 0;
      verilogPut_Key_1009 <= 0;
      verilogPut_FoundKey_1010 <= 0;
      verilogPut_Data_1011 <= 0;
      verilogPut_BtreeIndex_1012 <= 0;
      verilogPut_StuckIndex_1013 <= 0;
      verilogPut_MergeSuccess_1014 <= 0;
      verilogPut_childKey_1015 <= 0;
      verilogPut_size_1016 <= 0;
      verilogPut_childData_1017 <= 0;
      verilogPut_indexLeft_1018 <= 0;
      verilogPut_indexRight_1019 <= 0;
      verilogPut_midKey_1020 <= 0;
      verilogPut_success_1021 <= 0;
      verilogPut_test_1022 <= 0;
      verilogPut_next_1023 <= 0;
      verilogPut_root_1024 <= 0;
      verilogPut_isFree_1025 <= 0;
      verilogPut_index_1026 <= 0;
      verilogPut_size_1027 <= 0;
      verilogPut_isLeaf_1028 <= 0;
      verilogPut_nextFree_1029 <= 0;
      verilogPut_Key_0_1030 <= 0;
      verilogPut_KeyCompares_0_1031 <= 0;
      verilogPut_KeyCollapse_0_1032 <= 0;
      verilogPut_Data_0_1033 <= 0;
      verilogPut_Key_1_1034 <= 0;
      verilogPut_KeyCompares_1_1035 <= 0;
      verilogPut_KeyCollapse_1_1036 <= 0;
      verilogPut_Data_1_1037 <= 0;
      verilogPut_Key_2_1038 <= 0;
      verilogPut_KeyCompares_2_1039 <= 0;
      verilogPut_KeyCollapse_2_1040 <= 0;
      verilogPut_Data_2_1041 <= 0;
      verilogPut_Key_3_1042 <= 0;
      verilogPut_KeyCompares_3_1043 <= 0;
      verilogPut_KeyCollapse_3_1044 <= 0;
      verilogPut_Data_3_1045 <= 0;
      verilogPut_Found_1046 <= 0;
      verilogPut_Key_1047 <= 0;
      verilogPut_FoundKey_1048 <= 0;
      verilogPut_Data_1049 <= 0;
      verilogPut_BtreeIndex_1050 <= 0;
      verilogPut_StuckIndex_1051 <= 0;
      verilogPut_MergeSuccess_1052 <= 0;
      verilogPut_index_1053 <= 0;
      verilogPut_size_1054 <= 0;
      verilogPut_isLeaf_1055 <= 0;
      verilogPut_nextFree_1056 <= 0;
      verilogPut_Key_0_1057 <= 0;
      verilogPut_KeyCompares_0_1058 <= 0;
      verilogPut_KeyCollapse_0_1059 <= 0;
      verilogPut_Data_0_1060 <= 0;
      verilogPut_Key_1_1061 <= 0;
      verilogPut_KeyCompares_1_1062 <= 0;
      verilogPut_KeyCollapse_1_1063 <= 0;
      verilogPut_Data_1_1064 <= 0;
      verilogPut_Key_2_1065 <= 0;
      verilogPut_KeyCompares_2_1066 <= 0;
      verilogPut_KeyCollapse_2_1067 <= 0;
      verilogPut_Data_2_1068 <= 0;
      verilogPut_Key_3_1069 <= 0;
      verilogPut_KeyCompares_3_1070 <= 0;
      verilogPut_KeyCollapse_3_1071 <= 0;
      verilogPut_Data_3_1072 <= 0;
      verilogPut_Found_1073 <= 0;
      verilogPut_Key_1074 <= 0;
      verilogPut_FoundKey_1075 <= 0;
      verilogPut_Data_1076 <= 0;
      verilogPut_BtreeIndex_1077 <= 0;
      verilogPut_StuckIndex_1078 <= 0;
      verilogPut_MergeSuccess_1079 <= 0;
      verilogPut_childKey_1080 <= 0;
      verilogPut_size_1081 <= 0;
      verilogPut_childData_1082 <= 0;
      verilogPut_indexLeft_1083 <= 0;
      verilogPut_indexRight_1084 <= 0;
      verilogPut_midKey_1085 <= 0;
      verilogPut_success_1086 <= 0;
      verilogPut_test_1087 <= 0;
      verilogPut_next_1088 <= 0;
      verilogPut_root_1089 <= 0;
      verilogPut_isFree_1090 <= 0;
      verilogPut_index_1091 <= 0;
      verilogPut_size_1092 <= 0;
      verilogPut_isLeaf_1093 <= 0;
      verilogPut_nextFree_1094 <= 0;
      verilogPut_Key_0_1095 <= 0;
      verilogPut_KeyCompares_0_1096 <= 0;
      verilogPut_KeyCollapse_0_1097 <= 0;
      verilogPut_Data_0_1098 <= 0;
      verilogPut_Key_1_1099 <= 0;
      verilogPut_KeyCompares_1_1100 <= 0;
      verilogPut_KeyCollapse_1_1101 <= 0;
      verilogPut_Data_1_1102 <= 0;
      verilogPut_Key_2_1103 <= 0;
      verilogPut_KeyCompares_2_1104 <= 0;
      verilogPut_KeyCollapse_2_1105 <= 0;
      verilogPut_Data_2_1106 <= 0;
      verilogPut_Key_3_1107 <= 0;
      verilogPut_KeyCompares_3_1108 <= 0;
      verilogPut_KeyCollapse_3_1109 <= 0;
      verilogPut_Data_3_1110 <= 0;
      verilogPut_Found_1111 <= 0;
      verilogPut_Key_1112 <= 0;
      verilogPut_FoundKey_1113 <= 0;
      verilogPut_Data_1114 <= 0;
      verilogPut_BtreeIndex_1115 <= 0;
      verilogPut_StuckIndex_1116 <= 0;
      verilogPut_MergeSuccess_1117 <= 0;
      verilogPut_index_1118 <= 0;
      verilogPut_size_1119 <= 0;
      verilogPut_isLeaf_1120 <= 0;
      verilogPut_nextFree_1121 <= 0;
      verilogPut_Key_0_1122 <= 0;
      verilogPut_KeyCompares_0_1123 <= 0;
      verilogPut_KeyCollapse_0_1124 <= 0;
      verilogPut_Data_0_1125 <= 0;
      verilogPut_Key_1_1126 <= 0;
      verilogPut_KeyCompares_1_1127 <= 0;
      verilogPut_KeyCollapse_1_1128 <= 0;
      verilogPut_Data_1_1129 <= 0;
      verilogPut_Key_2_1130 <= 0;
      verilogPut_KeyCompares_2_1131 <= 0;
      verilogPut_KeyCollapse_2_1132 <= 0;
      verilogPut_Data_2_1133 <= 0;
      verilogPut_Key_3_1134 <= 0;
      verilogPut_KeyCompares_3_1135 <= 0;
      verilogPut_KeyCollapse_3_1136 <= 0;
      verilogPut_Data_3_1137 <= 0;
      verilogPut_Found_1138 <= 0;
      verilogPut_Key_1139 <= 0;
      verilogPut_FoundKey_1140 <= 0;
      verilogPut_Data_1141 <= 0;
      verilogPut_BtreeIndex_1142 <= 0;
      verilogPut_StuckIndex_1143 <= 0;
      verilogPut_MergeSuccess_1144 <= 0;
      verilogPut_childKey_1145 <= 0;
      verilogPut_childData_1146 <= 0;
      verilogPut_indexLeft_1147 <= 0;
      verilogPut_indexRight_1148 <= 0;
      verilogPut_midKey_1149 <= 0;
      verilogPut_success_1150 <= 0;
      verilogPut_test_1151 <= 0;
      verilogPut_next_1152 <= 0;
      verilogPut_root_1153 <= 0;
      verilogPut_isFree_1154 <= 0;
      verilogPut_index_1155 <= 0;
      verilogPut_size_1156 <= 0;
      verilogPut_isLeaf_1157 <= 0;
      verilogPut_nextFree_1158 <= 0;
      verilogPut_Key_0_1159 <= 0;
      verilogPut_KeyCompares_0_1160 <= 0;
      verilogPut_KeyCollapse_0_1161 <= 0;
      verilogPut_Data_0_1162 <= 0;
      verilogPut_Key_1_1163 <= 0;
      verilogPut_KeyCompares_1_1164 <= 0;
      verilogPut_KeyCollapse_1_1165 <= 0;
      verilogPut_Data_1_1166 <= 0;
      verilogPut_Key_2_1167 <= 0;
      verilogPut_KeyCompares_2_1168 <= 0;
      verilogPut_KeyCollapse_2_1169 <= 0;
      verilogPut_Data_2_1170 <= 0;
      verilogPut_Key_3_1171 <= 0;
      verilogPut_KeyCompares_3_1172 <= 0;
      verilogPut_KeyCollapse_3_1173 <= 0;
      verilogPut_Data_3_1174 <= 0;
      verilogPut_Found_1175 <= 0;
      verilogPut_Key_1176 <= 0;
      verilogPut_FoundKey_1177 <= 0;
      verilogPut_Data_1178 <= 0;
      verilogPut_BtreeIndex_1179 <= 0;
      verilogPut_StuckIndex_1180 <= 0;
      verilogPut_MergeSuccess_1181 <= 0;
      verilogPut_index_1182 <= 0;
      verilogPut_size_1183 <= 0;
      verilogPut_isLeaf_1184 <= 0;
      verilogPut_nextFree_1185 <= 0;
      verilogPut_Key_0_1186 <= 0;
      verilogPut_KeyCompares_0_1187 <= 0;
      verilogPut_KeyCollapse_0_1188 <= 0;
      verilogPut_Data_0_1189 <= 0;
      verilogPut_Key_1_1190 <= 0;
      verilogPut_KeyCompares_1_1191 <= 0;
      verilogPut_KeyCollapse_1_1192 <= 0;
      verilogPut_Data_1_1193 <= 0;
      verilogPut_Key_2_1194 <= 0;
      verilogPut_KeyCompares_2_1195 <= 0;
      verilogPut_KeyCollapse_2_1196 <= 0;
      verilogPut_Data_2_1197 <= 0;
      verilogPut_Key_3_1198 <= 0;
      verilogPut_KeyCompares_3_1199 <= 0;
      verilogPut_KeyCollapse_3_1200 <= 0;
      verilogPut_Data_3_1201 <= 0;
      verilogPut_Found_1202 <= 0;
      verilogPut_Key_1203 <= 0;
      verilogPut_FoundKey_1204 <= 0;
      verilogPut_Data_1205 <= 0;
      verilogPut_BtreeIndex_1206 <= 0;
      verilogPut_StuckIndex_1207 <= 0;
      verilogPut_MergeSuccess_1208 <= 0;
      verilogPut_childKey_1209 <= 0;
      verilogPut_leftChild_1210 <= 0;
      verilogPut_rightChild_1211 <= 0;
      verilogPut_childData_1212 <= 0;
      verilogPut_indexLeft_1213 <= 0;
      verilogPut_indexRight_1214 <= 0;
      verilogPut_midKey_1215 <= 0;
      verilogPut_success_1216 <= 0;
      verilogPut_test_1217 <= 0;
      verilogPut_next_1218 <= 0;
      verilogPut_root_1219 <= 0;
      verilogPut_isFree_1220 <= 0;
      verilogPut_index_1221 <= 0;
      verilogPut_size_1222 <= 0;
      verilogPut_isLeaf_1223 <= 0;
      verilogPut_nextFree_1224 <= 0;
      verilogPut_Key_0_1225 <= 0;
      verilogPut_KeyCompares_0_1226 <= 0;
      verilogPut_KeyCollapse_0_1227 <= 0;
      verilogPut_Data_0_1228 <= 0;
      verilogPut_Key_1_1229 <= 0;
      verilogPut_KeyCompares_1_1230 <= 0;
      verilogPut_KeyCollapse_1_1231 <= 0;
      verilogPut_Data_1_1232 <= 0;
      verilogPut_Key_2_1233 <= 0;
      verilogPut_KeyCompares_2_1234 <= 0;
      verilogPut_KeyCollapse_2_1235 <= 0;
      verilogPut_Data_2_1236 <= 0;
      verilogPut_Key_3_1237 <= 0;
      verilogPut_KeyCompares_3_1238 <= 0;
      verilogPut_KeyCollapse_3_1239 <= 0;
      verilogPut_Data_3_1240 <= 0;
      verilogPut_Found_1241 <= 0;
      verilogPut_Key_1242 <= 0;
      verilogPut_FoundKey_1243 <= 0;
      verilogPut_Data_1244 <= 0;
      verilogPut_BtreeIndex_1245 <= 0;
      verilogPut_StuckIndex_1246 <= 0;
      verilogPut_MergeSuccess_1247 <= 0;
      verilogPut_index_1248 <= 0;
      verilogPut_size_1249 <= 0;
      verilogPut_isLeaf_1250 <= 0;
      verilogPut_nextFree_1251 <= 0;
      verilogPut_Key_0_1252 <= 0;
      verilogPut_KeyCompares_0_1253 <= 0;
      verilogPut_KeyCollapse_0_1254 <= 0;
      verilogPut_Data_0_1255 <= 0;
      verilogPut_Key_1_1256 <= 0;
      verilogPut_KeyCompares_1_1257 <= 0;
      verilogPut_KeyCollapse_1_1258 <= 0;
      verilogPut_Data_1_1259 <= 0;
      verilogPut_Key_2_1260 <= 0;
      verilogPut_KeyCompares_2_1261 <= 0;
      verilogPut_KeyCollapse_2_1262 <= 0;
      verilogPut_Data_2_1263 <= 0;
      verilogPut_Key_3_1264 <= 0;
      verilogPut_KeyCompares_3_1265 <= 0;
      verilogPut_KeyCollapse_3_1266 <= 0;
      verilogPut_Data_3_1267 <= 0;
      verilogPut_Found_1268 <= 0;
      verilogPut_Key_1269 <= 0;
      verilogPut_FoundKey_1270 <= 0;
      verilogPut_Data_1271 <= 0;
      verilogPut_BtreeIndex_1272 <= 0;
      verilogPut_StuckIndex_1273 <= 0;
      verilogPut_MergeSuccess_1274 <= 0;
      verilogPut_childKey_1275 <= 0;
      verilogPut_childData_1276 <= 0;
      verilogPut_indexLeft_1277 <= 0;
      verilogPut_indexRight_1278 <= 0;
      verilogPut_midKey_1279 <= 0;
      verilogPut_success_1280 <= 0;
      verilogPut_test_1281 <= 0;
      verilogPut_next_1282 <= 0;
      verilogPut_root_1283 <= 0;
      verilogPut_isFree_1284 <= 0;
      verilogPut_index_1285 <= 0;
      verilogPut_size_1286 <= 0;
      verilogPut_isLeaf_1287 <= 0;
      verilogPut_nextFree_1288 <= 0;
      verilogPut_Key_0_1289 <= 0;
      verilogPut_KeyCompares_0_1290 <= 0;
      verilogPut_KeyCollapse_0_1291 <= 0;
      verilogPut_Data_0_1292 <= 0;
      verilogPut_Key_1_1293 <= 0;
      verilogPut_KeyCompares_1_1294 <= 0;
      verilogPut_KeyCollapse_1_1295 <= 0;
      verilogPut_Data_1_1296 <= 0;
      verilogPut_Key_2_1297 <= 0;
      verilogPut_KeyCompares_2_1298 <= 0;
      verilogPut_KeyCollapse_2_1299 <= 0;
      verilogPut_Data_2_1300 <= 0;
      verilogPut_Key_3_1301 <= 0;
      verilogPut_KeyCompares_3_1302 <= 0;
      verilogPut_KeyCollapse_3_1303 <= 0;
      verilogPut_Data_3_1304 <= 0;
      verilogPut_Found_1305 <= 0;
      verilogPut_Key_1306 <= 0;
      verilogPut_FoundKey_1307 <= 0;
      verilogPut_Data_1308 <= 0;
      verilogPut_BtreeIndex_1309 <= 0;
      verilogPut_StuckIndex_1310 <= 0;
      verilogPut_MergeSuccess_1311 <= 0;
      verilogPut_index_1312 <= 0;
      verilogPut_size_1313 <= 0;
      verilogPut_isLeaf_1314 <= 0;
      verilogPut_nextFree_1315 <= 0;
      verilogPut_Key_0_1316 <= 0;
      verilogPut_KeyCompares_0_1317 <= 0;
      verilogPut_KeyCollapse_0_1318 <= 0;
      verilogPut_Data_0_1319 <= 0;
      verilogPut_Key_1_1320 <= 0;
      verilogPut_KeyCompares_1_1321 <= 0;
      verilogPut_KeyCollapse_1_1322 <= 0;
      verilogPut_Data_1_1323 <= 0;
      verilogPut_Key_2_1324 <= 0;
      verilogPut_KeyCompares_2_1325 <= 0;
      verilogPut_KeyCollapse_2_1326 <= 0;
      verilogPut_Data_2_1327 <= 0;
      verilogPut_Key_3_1328 <= 0;
      verilogPut_KeyCompares_3_1329 <= 0;
      verilogPut_KeyCollapse_3_1330 <= 0;
      verilogPut_Data_3_1331 <= 0;
      verilogPut_Found_1332 <= 0;
      verilogPut_Key_1333 <= 0;
      verilogPut_FoundKey_1334 <= 0;
      verilogPut_Data_1335 <= 0;
      verilogPut_BtreeIndex_1336 <= 0;
      verilogPut_StuckIndex_1337 <= 0;
      verilogPut_MergeSuccess_1338 <= 0;
      verilogPut_childKey_1339 <= 0;
      verilogPut_leftChild_1340 <= 0;
      verilogPut_rightChild_1341 <= 0;
      verilogPut_childData_1342 <= 0;
      verilogPut_indexLeft_1343 <= 0;
      verilogPut_indexRight_1344 <= 0;
      verilogPut_midKey_1345 <= 0;
      verilogPut_success_1346 <= 0;
      verilogPut_test_1347 <= 0;
      verilogPut_next_1348 <= 0;
      verilogPut_root_1349 <= 0;
      verilogPut_isFree_1350 <= 0;
      verilogPut_index_1351 <= 0;
      verilogPut_size_1352 <= 0;
      verilogPut_isLeaf_1353 <= 0;
      verilogPut_nextFree_1354 <= 0;
      verilogPut_Key_0_1355 <= 0;
      verilogPut_KeyCompares_0_1356 <= 0;
      verilogPut_KeyCollapse_0_1357 <= 0;
      verilogPut_Data_0_1358 <= 0;
      verilogPut_Key_1_1359 <= 0;
      verilogPut_KeyCompares_1_1360 <= 0;
      verilogPut_KeyCollapse_1_1361 <= 0;
      verilogPut_Data_1_1362 <= 0;
      verilogPut_Key_2_1363 <= 0;
      verilogPut_KeyCompares_2_1364 <= 0;
      verilogPut_KeyCollapse_2_1365 <= 0;
      verilogPut_Data_2_1366 <= 0;
      verilogPut_Key_3_1367 <= 0;
      verilogPut_KeyCompares_3_1368 <= 0;
      verilogPut_KeyCollapse_3_1369 <= 0;
      verilogPut_Data_3_1370 <= 0;
      verilogPut_Found_1371 <= 0;
      verilogPut_Key_1372 <= 0;
      verilogPut_FoundKey_1373 <= 0;
      verilogPut_Data_1374 <= 0;
      verilogPut_BtreeIndex_1375 <= 0;
      verilogPut_StuckIndex_1376 <= 0;
      verilogPut_MergeSuccess_1377 <= 0;
      verilogPut_index_1378 <= 0;
      verilogPut_size_1379 <= 0;
      verilogPut_isLeaf_1380 <= 0;
      verilogPut_nextFree_1381 <= 0;
      verilogPut_Key_0_1382 <= 0;
      verilogPut_KeyCompares_0_1383 <= 0;
      verilogPut_KeyCollapse_0_1384 <= 0;
      verilogPut_Data_0_1385 <= 0;
      verilogPut_Key_1_1386 <= 0;
      verilogPut_KeyCompares_1_1387 <= 0;
      verilogPut_KeyCollapse_1_1388 <= 0;
      verilogPut_Data_1_1389 <= 0;
      verilogPut_Key_2_1390 <= 0;
      verilogPut_KeyCompares_2_1391 <= 0;
      verilogPut_KeyCollapse_2_1392 <= 0;
      verilogPut_Data_2_1393 <= 0;
      verilogPut_Key_3_1394 <= 0;
      verilogPut_KeyCompares_3_1395 <= 0;
      verilogPut_KeyCollapse_3_1396 <= 0;
      verilogPut_Data_3_1397 <= 0;
      verilogPut_Found_1398 <= 0;
      verilogPut_Key_1399 <= 0;
      verilogPut_FoundKey_1400 <= 0;
      verilogPut_Data_1401 <= 0;
      verilogPut_BtreeIndex_1402 <= 0;
      verilogPut_StuckIndex_1403 <= 0;
      verilogPut_MergeSuccess_1404 <= 0;
      verilogPut_childKey_1405 <= 0;
      verilogPut_childData_1406 <= 0;
      verilogPut_indexLeft_1407 <= 0;
      verilogPut_indexRight_1408 <= 0;
      verilogPut_midKey_1409 <= 0;
      verilogPut_success_1410 <= 0;
      verilogPut_test_1411 <= 0;
      verilogPut_next_1412 <= 0;
      verilogPut_root_1413 <= 0;
      verilogPut_isFree_1414 <= 0;
      verilogPut_index_1415 <= 0;
      verilogPut_size_1416 <= 0;
      verilogPut_isLeaf_1417 <= 0;
      verilogPut_nextFree_1418 <= 0;
      verilogPut_Key_0_1419 <= 0;
      verilogPut_KeyCompares_0_1420 <= 0;
      verilogPut_KeyCollapse_0_1421 <= 0;
      verilogPut_Data_0_1422 <= 0;
      verilogPut_Key_1_1423 <= 0;
      verilogPut_KeyCompares_1_1424 <= 0;
      verilogPut_KeyCollapse_1_1425 <= 0;
      verilogPut_Data_1_1426 <= 0;
      verilogPut_Key_2_1427 <= 0;
      verilogPut_KeyCompares_2_1428 <= 0;
      verilogPut_KeyCollapse_2_1429 <= 0;
      verilogPut_Data_2_1430 <= 0;
      verilogPut_Key_3_1431 <= 0;
      verilogPut_KeyCompares_3_1432 <= 0;
      verilogPut_KeyCollapse_3_1433 <= 0;
      verilogPut_Data_3_1434 <= 0;
      verilogPut_Found_1435 <= 0;
      verilogPut_Key_1436 <= 0;
      verilogPut_FoundKey_1437 <= 0;
      verilogPut_Data_1438 <= 0;
      verilogPut_BtreeIndex_1439 <= 0;
      verilogPut_StuckIndex_1440 <= 0;
      verilogPut_MergeSuccess_1441 <= 0;
      verilogPut_index_1442 <= 0;
      verilogPut_size_1443 <= 0;
      verilogPut_isLeaf_1444 <= 0;
      verilogPut_nextFree_1445 <= 0;
      verilogPut_Key_0_1446 <= 0;
      verilogPut_KeyCompares_0_1447 <= 0;
      verilogPut_KeyCollapse_0_1448 <= 0;
      verilogPut_Data_0_1449 <= 0;
      verilogPut_Key_1_1450 <= 0;
      verilogPut_KeyCompares_1_1451 <= 0;
      verilogPut_KeyCollapse_1_1452 <= 0;
      verilogPut_Data_1_1453 <= 0;
      verilogPut_Key_2_1454 <= 0;
      verilogPut_KeyCompares_2_1455 <= 0;
      verilogPut_KeyCollapse_2_1456 <= 0;
      verilogPut_Data_2_1457 <= 0;
      verilogPut_Key_3_1458 <= 0;
      verilogPut_KeyCompares_3_1459 <= 0;
      verilogPut_KeyCollapse_3_1460 <= 0;
      verilogPut_Data_3_1461 <= 0;
      verilogPut_Found_1462 <= 0;
      verilogPut_Key_1463 <= 0;
      verilogPut_FoundKey_1464 <= 0;
      verilogPut_Data_1465 <= 0;
      verilogPut_BtreeIndex_1466 <= 0;
      verilogPut_StuckIndex_1467 <= 0;
      verilogPut_MergeSuccess_1468 <= 0;
      verilogPut_childKey_1469 <= 0;
      verilogPut_leftChild_1470 <= 0;
      verilogPut_rightChild_1471 <= 0;
      verilogPut_childData_1472 <= 0;
      verilogPut_indexLeft_1473 <= 0;
      verilogPut_indexRight_1474 <= 0;
      verilogPut_midKey_1475 <= 0;
      verilogPut_success_1476 <= 0;
      verilogPut_test_1477 <= 0;
      verilogPut_next_1478 <= 0;
      verilogPut_root_1479 <= 0;
      verilogPut_isFree_1480 <= 0;
      stuckIsLeaf_7_requestedAt <= -1;
      stuckIsLeaf_8_requestedAt <= -1;
      stuckIsFree_11_requestedAt <= -1;
      freeNext_9_requestedAt <= -1;
      freeNext_10_requestedAt <= -1;
      stuckSize_5_requestedAt <= -1;
      stuckSize_6_requestedAt <= -1;
      stuckKeys_1_requestedAt <= -1;
      stuckKeys_2_requestedAt <= -1;
      stuckData_3_requestedAt <= -1;
      stuckData_4_requestedAt <= -1;
    end
    else begin                                   // Run the process in full parallel
      case(verilogPut_pc)
        0: begin
          verilogPut_k_0 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        1: begin
          verilogPut_d_1 <= 11;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        2: begin
          verilogPut_BtreeIndex_98 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        3: begin
          verilogPut_index_74 <= verilogPut_BtreeIndex_98;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        4: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_74;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_74;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_74;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_74;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        5: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        6: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        7: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        8: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        9: begin
          verilogPut_size_75 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_76 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_78 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_81 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_82 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_85 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_86 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_89 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_90 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_93 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        10: begin
          if (verilogPut_isLeaf_76 == 0) begin
            verilogPut_pc <= 17;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        11: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 == verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 == verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 == verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 == verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        12: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        13: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        14: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Key_95 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Key_95 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Key_95 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Key_95 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        15: begin
          verilogPut_pc <= 23;
        end
        16: begin
          verilogPut_pc <= 23;
        end
        17: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 <= verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 >  verilogPut_Key_0_78 && verilogPut_k_0 <= verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 >  verilogPut_Key_1_82 && verilogPut_k_0 <= verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 >  verilogPut_Key_2_86 && verilogPut_k_0 <= verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        18: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        19: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        20: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_FoundKey_96 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_FoundKey_96 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_FoundKey_96 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_FoundKey_96 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
            case (verilogPut_size_75)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        21: begin
          verilogPut_BtreeIndex_98 <= verilogPut_Data_97;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        22: begin
          verilogPut_pc <= 3;
        end
        23: begin
          if (verilogPut_Found_94 == 0) begin
            verilogPut_pc <= 26;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        24: begin
          if (verilogPut_StuckIndex_99 == verilogPut_size_75) begin
            verilogPut_size_75 <= verilogPut_size_75+1;
          end
          case (verilogPut_StuckIndex_99)
            0: begin
              verilogPut_Key_0_78 <= verilogPut_k_0;
              verilogPut_Data_0_81 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_82 <= verilogPut_k_0;
              verilogPut_Data_1_85 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_86 <= verilogPut_k_0;
              verilogPut_Data_2_89 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_90 <= verilogPut_k_0;
              verilogPut_Data_3_93 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        25: begin
          verilogPut_pc <= 37;
        end
        26: begin
          verilogPut_notFull_107 <= verilogPut_size_75< 4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        27: begin
          if (verilogPut_notFull_107 == 0) begin
            verilogPut_pc <= 36;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        28: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 <= verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 >  verilogPut_Key_0_78 && verilogPut_k_0 <= verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 >  verilogPut_Key_1_82 && verilogPut_k_0 <= verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 >  verilogPut_Key_2_86 && verilogPut_k_0 <= verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        29: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        30: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        31: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_FoundKey_96 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_FoundKey_96 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_FoundKey_96 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_FoundKey_96 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
            case (verilogPut_size_75)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        32: begin
          verilogPut_size_75 <= verilogPut_size_75+1;
          if (3 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_3_90 <= verilogPut_Key_2_86;
            verilogPut_Data_3_93 <= verilogPut_Data_2_89;
          end
          if (2 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_2_86 <= verilogPut_Key_1_82;
            verilogPut_Data_2_89 <= verilogPut_Data_1_85;
          end
          if (1 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_1_82 <= verilogPut_Key_0_78;
            verilogPut_Data_1_85 <= verilogPut_Data_0_81;
          end
          case (verilogPut_StuckIndex_99)
            0: begin
              verilogPut_Key_0_78 <= verilogPut_k_0;
              verilogPut_Data_0_81 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_82 <= verilogPut_k_0;
              verilogPut_Data_1_85 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_86 <= verilogPut_k_0;
              verilogPut_Data_2_89 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_90 <= verilogPut_k_0;
              verilogPut_Data_3_93 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        33: begin
          verilogPut_Found_94 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        34: begin
          verilogPut_pc <= verilogPut_pc + 1;
        end
        35: begin
          verilogPut_pc <= 37;
        end
        36: begin
          verilogPut_pc <= 41;
        end
        37: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_74;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_75;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_74;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_78;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_82;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_86;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_90;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_74;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_81;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_85;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_89;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_93;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        38: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        39: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        40: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        41: begin
          if (verilogPut_Found_94 >  0) begin
            verilogPut_pc <= 449;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        42: begin
          if (verilogPut_BtreeIndex_98 == 0) begin
            verilogPut_pc <= 44;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        43: begin
          verilogPut_pc <= 137;
        end
        44: begin
          verilogPut_index_108 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        45: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_108;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_108;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_108;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_108;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        46: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        47: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        48: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        49: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        50: begin
          verilogPut_size_109 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_110 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_112 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_115 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_116 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_119 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_120 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_123 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_124 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_127 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        51: begin
          if (verilogPut_size_109 < 4) begin
            verilogPut_pc <= 97;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        52: begin
          verilogPut_Key_0_139 <= verilogPut_Key_0_112;
          verilogPut_Data_0_142 <= verilogPut_Data_0_115;
          verilogPut_Key_1_143 <= verilogPut_Key_1_116;
          verilogPut_Data_1_146 <= verilogPut_Data_1_119;
          verilogPut_size_136 <= 2;
          verilogPut_Key_0_166 <= verilogPut_Key_2_120;
          verilogPut_Data_0_169 <= verilogPut_Data_2_123;
          verilogPut_Key_1_170 <= verilogPut_Key_3_124;
          verilogPut_Data_1_173 <= verilogPut_Data_3_127;
          verilogPut_size_163 <= 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        53: begin
          verilogPut_root_197 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        54: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_197;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        55: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        56: begin
          verilogPut_indexLeft_189 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        57: begin
          if (verilogPut_indexLeft_189 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_199 <= 1;
          verilogPut_isFree_200 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        58: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexLeft_189;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexLeft_189;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_199;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_189;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_200;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        59: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        60: begin
          verilogPut_next_198 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        61: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_197;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_198;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        62: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        63: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        64: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        65: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexLeft_189;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_136;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexLeft_189;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_139;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_143;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_147;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_151;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexLeft_189;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_142;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_146;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_150;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_154;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        66: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        67: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        68: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        69: begin
          verilogPut_root_201 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        70: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_201;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        71: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        72: begin
          verilogPut_indexRight_190 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        73: begin
          if (verilogPut_indexRight_190 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_203 <= 1;
          verilogPut_isFree_204 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        74: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexRight_190;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexRight_190;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_203;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_190;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_204;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        75: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        76: begin
          verilogPut_next_202 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        77: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_201;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_202;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        78: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        79: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        80: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        81: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexRight_190;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_163;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexRight_190;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_166;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_170;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_174;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_178;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexRight_190;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_169;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_173;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_177;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_181;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        82: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        83: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        84: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        85: begin
          case (verilogPut_size_136)
            1: begin
              verilogPut_Key_156 <= verilogPut_Key_0_139;
              verilogPut_Data_158 <= verilogPut_Data_0_142;
            end
            2: begin
              verilogPut_Key_156 <= verilogPut_Key_1_143;
              verilogPut_Data_158 <= verilogPut_Data_1_146;
            end
            3: begin
              verilogPut_Key_156 <= verilogPut_Key_2_147;
              verilogPut_Data_158 <= verilogPut_Data_2_150;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        86: begin
          verilogPut_Key_183 <= verilogPut_Key_0_166;
          verilogPut_Data_185 <= verilogPut_Data_0_169;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        87: begin
          verilogPut_midKey_191 <= (verilogPut_Key_156 + verilogPut_Key_183) / 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        88: begin
          verilogPut_size_109 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        89: begin
          case (verilogPut_size_109)
            0: begin
              verilogPut_Key_0_112 <= verilogPut_midKey_191;
              verilogPut_Data_0_115 <= verilogPut_indexLeft_189;
            end
            1: begin
              verilogPut_Key_1_116 <= verilogPut_midKey_191;
              verilogPut_Data_1_119 <= verilogPut_indexLeft_189;
            end
            2: begin
              verilogPut_Key_2_120 <= verilogPut_midKey_191;
              verilogPut_Data_2_123 <= verilogPut_indexLeft_189;
            end
            3: begin
              verilogPut_Key_3_124 <= verilogPut_midKey_191;
              verilogPut_Data_3_127 <= verilogPut_indexLeft_189;
            end
          endcase
          verilogPut_size_109 <= verilogPut_size_109+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        90: begin
          case (verilogPut_size_109)
            0: begin
              verilogPut_Key_0_112 <= verilogPut_midKey_191;
              verilogPut_Data_0_115 <= verilogPut_indexRight_190;
            end
            1: begin
              verilogPut_Key_1_116 <= verilogPut_midKey_191;
              verilogPut_Data_1_119 <= verilogPut_indexRight_190;
            end
            2: begin
              verilogPut_Key_2_120 <= verilogPut_midKey_191;
              verilogPut_Data_2_123 <= verilogPut_indexRight_190;
            end
            3: begin
              verilogPut_Key_3_124 <= verilogPut_midKey_191;
              verilogPut_Data_3_127 <= verilogPut_indexRight_190;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        91: begin
          verilogPut_isLeaf_110 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        92: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_108;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_109;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_index_108;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_110;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_108;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_112;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_116;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_120;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_124;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_108;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_115;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_119;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_123;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_127;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        93: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        94: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        95: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        96: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        97: begin
          verilogPut_BtreeIndex_98 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        98: begin
          verilogPut_index_74 <= verilogPut_BtreeIndex_98;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        99: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_74;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_74;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_74;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_74;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        100: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        101: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        102: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        103: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        104: begin
          verilogPut_size_75 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_76 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_78 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_81 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_82 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_85 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_86 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_89 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_90 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_93 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        105: begin
          if (verilogPut_isLeaf_76 == 0) begin
            verilogPut_pc <= 112;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        106: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 == verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 == verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 == verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 == verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        107: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        108: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        109: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Key_95 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Key_95 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Key_95 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Key_95 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        110: begin
          verilogPut_pc <= 118;
        end
        111: begin
          verilogPut_pc <= 118;
        end
        112: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 <= verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 >  verilogPut_Key_0_78 && verilogPut_k_0 <= verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 >  verilogPut_Key_1_82 && verilogPut_k_0 <= verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 >  verilogPut_Key_2_86 && verilogPut_k_0 <= verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        113: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        114: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        115: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_FoundKey_96 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_FoundKey_96 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_FoundKey_96 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_FoundKey_96 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
            case (verilogPut_size_75)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        116: begin
          verilogPut_BtreeIndex_98 <= verilogPut_Data_97;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        117: begin
          verilogPut_pc <= 98;
        end
        118: begin
          if (verilogPut_Found_94 == 0) begin
            verilogPut_pc <= 121;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        119: begin
          if (verilogPut_StuckIndex_99 == verilogPut_size_75) begin
            verilogPut_size_75 <= verilogPut_size_75+1;
          end
          case (verilogPut_StuckIndex_99)
            0: begin
              verilogPut_Key_0_78 <= verilogPut_k_0;
              verilogPut_Data_0_81 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_82 <= verilogPut_k_0;
              verilogPut_Data_1_85 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_86 <= verilogPut_k_0;
              verilogPut_Data_2_89 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_90 <= verilogPut_k_0;
              verilogPut_Data_3_93 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        120: begin
          verilogPut_pc <= 132;
        end
        121: begin
          verilogPut_notFull_206 <= verilogPut_size_75< 4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        122: begin
          if (verilogPut_notFull_206 == 0) begin
            verilogPut_pc <= 131;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        123: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 <= verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 >  verilogPut_Key_0_78 && verilogPut_k_0 <= verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 >  verilogPut_Key_1_82 && verilogPut_k_0 <= verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 >  verilogPut_Key_2_86 && verilogPut_k_0 <= verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        124: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        125: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        126: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_FoundKey_96 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_FoundKey_96 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_FoundKey_96 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_FoundKey_96 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
            case (verilogPut_size_75)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        127: begin
          verilogPut_size_75 <= verilogPut_size_75+1;
          if (3 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_3_90 <= verilogPut_Key_2_86;
            verilogPut_Data_3_93 <= verilogPut_Data_2_89;
          end
          if (2 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_2_86 <= verilogPut_Key_1_82;
            verilogPut_Data_2_89 <= verilogPut_Data_1_85;
          end
          if (1 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_1_82 <= verilogPut_Key_0_78;
            verilogPut_Data_1_85 <= verilogPut_Data_0_81;
          end
          case (verilogPut_StuckIndex_99)
            0: begin
              verilogPut_Key_0_78 <= verilogPut_k_0;
              verilogPut_Data_0_81 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_82 <= verilogPut_k_0;
              verilogPut_Data_1_85 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_86 <= verilogPut_k_0;
              verilogPut_Data_2_89 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_90 <= verilogPut_k_0;
              verilogPut_Data_3_93 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        128: begin
          verilogPut_Found_94 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        129: begin
          verilogPut_pc <= verilogPut_pc + 1;
        end
        130: begin
          verilogPut_pc <= 132;
        end
        131: begin
          verilogPut_pc <= 136;
        end
        132: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_74;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_75;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_74;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_78;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_82;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_86;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_90;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_74;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_81;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_85;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_89;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_93;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        133: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        134: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        135: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        136: begin
          verilogPut_pc <= 449;
        end
        137: begin
          verilogPut_index_2 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        138: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_2;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_2;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_2;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_2;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        139: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        140: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        141: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        142: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        143: begin
          verilogPut_size_3 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_4 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_6 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_9 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_10 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_13 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_14 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_17 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_18 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_21 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        144: begin
          verilogPut_full_105 <= verilogPut_size_3>=3 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        145: begin
          if (verilogPut_full_105 == 0) begin
            verilogPut_pc <= 197;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        146: begin
          verilogPut_index_207 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        147: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_207;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_207;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_207;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_207;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        148: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        149: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        150: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        151: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        152: begin
          verilogPut_size_208 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_209 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_211 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_214 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_215 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_218 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_219 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_222 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_223 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_226 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        153: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        154: begin
          verilogPut_Key_0_238 <= verilogPut_Key_0_211;
          verilogPut_Data_0_241 <= verilogPut_Data_0_214;
          verilogPut_size_235 <= 1;
          verilogPut_Data_1_245 <= verilogPut_Data_1_218;
          verilogPut_Key_0_265 <= verilogPut_Key_2_219;
          verilogPut_Data_0_268 <= verilogPut_Data_2_222;
          case (verilogPut_size_208)
            0: begin
              verilogPut_size_262 <= -2;
              verilogPut_Data_1_272 <= verilogPut_Data_3_226;
            end
            1: begin
              verilogPut_size_262 <= -1;
              verilogPut_Data_1_272 <= verilogPut_Data_3_226;
            end
            2: begin
              verilogPut_size_262 <= 0;
              verilogPut_Data_1_272 <= verilogPut_Data_3_226;
            end
            3: begin
              verilogPut_size_262 <= 1;
              verilogPut_Data_1_272 <= verilogPut_Data_3_226;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        155: begin
          verilogPut_root_291 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        156: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_291;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        157: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        158: begin
          verilogPut_indexLeft_288 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        159: begin
          if (verilogPut_indexLeft_288 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_293 <= 0;
          verilogPut_isFree_294 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        160: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexLeft_288;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexLeft_288;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_293;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_288;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_294;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        161: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        162: begin
          verilogPut_next_292 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        163: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_291;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_292;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        164: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        165: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        166: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        167: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexLeft_288;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_235;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexLeft_288;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_238;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_242;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_246;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_250;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexLeft_288;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_241;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_245;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_249;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_253;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        168: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        169: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        170: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        171: begin
          verilogPut_root_295 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        172: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_295;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        173: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        174: begin
          verilogPut_indexRight_289 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        175: begin
          if (verilogPut_indexRight_289 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_297 <= 0;
          verilogPut_isFree_298 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        176: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexRight_289;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexRight_289;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_297;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_289;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_298;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        177: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        178: begin
          verilogPut_next_296 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        179: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_295;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_296;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        180: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        181: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        182: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        183: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexRight_289;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_262;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexRight_289;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_265;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_269;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_273;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_277;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexRight_289;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_268;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_272;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_276;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_280;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        184: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        185: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        186: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        187: begin
          verilogPut_midKey_290 <= verilogPut_Key_1_215;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        188: begin
          verilogPut_size_208 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        189: begin
          case (verilogPut_size_208)
            0: begin
              verilogPut_Key_0_211 <= verilogPut_midKey_290;
              verilogPut_Data_0_214 <= verilogPut_indexLeft_288;
            end
            1: begin
              verilogPut_Key_1_215 <= verilogPut_midKey_290;
              verilogPut_Data_1_218 <= verilogPut_indexLeft_288;
            end
            2: begin
              verilogPut_Key_2_219 <= verilogPut_midKey_290;
              verilogPut_Data_2_222 <= verilogPut_indexLeft_288;
            end
            3: begin
              verilogPut_Key_3_223 <= verilogPut_midKey_290;
              verilogPut_Data_3_226 <= verilogPut_indexLeft_288;
            end
          endcase
          verilogPut_size_208 <= verilogPut_size_208+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        190: begin
          case (verilogPut_size_208)
            0: begin
              verilogPut_Key_0_211 <= verilogPut_midKey_290;
              verilogPut_Data_0_214 <= verilogPut_indexRight_289;
            end
            1: begin
              verilogPut_Key_1_215 <= verilogPut_midKey_290;
              verilogPut_Data_1_218 <= verilogPut_indexRight_289;
            end
            2: begin
              verilogPut_Key_2_219 <= verilogPut_midKey_290;
              verilogPut_Data_2_222 <= verilogPut_indexRight_289;
            end
            3: begin
              verilogPut_Key_3_223 <= verilogPut_midKey_290;
              verilogPut_Data_3_226 <= verilogPut_indexRight_289;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        191: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_207;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_208;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_207;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_211;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_215;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_219;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_223;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_207;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_214;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_218;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_222;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_226;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        192: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        193: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        194: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        195: begin
          verilogPut_pc <= 41;
        end
        196: begin
          verilogPut_pc <= 197;
        end
        197: begin
          verilogPut_parent_102 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        198: begin
          verilogPut_index_2 <= verilogPut_parent_102;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        199: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_2;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_2;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_2;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_2;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        200: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        201: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        202: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        203: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        204: begin
          verilogPut_size_3 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_4 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_6 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_9 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_10 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_13 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_14 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_17 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_18 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_21 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        205: begin
          verilogPut_KeyCompares_0_7 <= verilogPut_k_0 <= verilogPut_Key_0_6 && 0 < verilogPut_size_3;
          verilogPut_KeyCollapse_0_8 <= 0;
          verilogPut_KeyCompares_1_11 <= verilogPut_k_0 >  verilogPut_Key_0_6 && verilogPut_k_0 <= verilogPut_Key_1_10 && 1 < verilogPut_size_3;
          verilogPut_KeyCollapse_1_12 <= 1;
          verilogPut_KeyCompares_2_15 <= verilogPut_k_0 >  verilogPut_Key_1_10 && verilogPut_k_0 <= verilogPut_Key_2_14 && 2 < verilogPut_size_3;
          verilogPut_KeyCollapse_2_16 <= 2;
          verilogPut_KeyCompares_3_19 <= verilogPut_k_0 >  verilogPut_Key_2_14 && verilogPut_k_0 <= verilogPut_Key_3_18 && 3 < verilogPut_size_3;
          verilogPut_KeyCollapse_3_20 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        206: begin
          if (verilogPut_KeyCompares_1_11) begin
            verilogPut_KeyCompares_0_7 <= 1;
            verilogPut_KeyCollapse_0_8 <= verilogPut_KeyCollapse_1_12;
          end
          if (verilogPut_KeyCompares_3_19) begin
            verilogPut_KeyCompares_2_15 <= 1;
            verilogPut_KeyCollapse_2_16 <= verilogPut_KeyCollapse_3_20;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        207: begin
          if (verilogPut_KeyCompares_2_15) begin
            verilogPut_KeyCompares_0_7 <= 1;
            verilogPut_KeyCollapse_0_8 <= verilogPut_KeyCollapse_2_16;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        208: begin
          if (verilogPut_KeyCompares_0_7) begin
            verilogPut_Found_40 <= 1;
            case (verilogPut_KeyCollapse_0_8)
              0: begin
                verilogPut_StuckIndex_45 <= 0;
                verilogPut_FoundKey_42 <= verilogPut_Key_0_6;
                verilogPut_Data_43 <= verilogPut_Data_0_9;
              end
              1: begin
                verilogPut_StuckIndex_45 <= 1;
                verilogPut_FoundKey_42 <= verilogPut_Key_1_10;
                verilogPut_Data_43 <= verilogPut_Data_1_13;
              end
              2: begin
                verilogPut_StuckIndex_45 <= 2;
                verilogPut_FoundKey_42 <= verilogPut_Key_2_14;
                verilogPut_Data_43 <= verilogPut_Data_2_17;
              end
              3: begin
                verilogPut_StuckIndex_45 <= 3;
                verilogPut_FoundKey_42 <= verilogPut_Key_3_18;
                verilogPut_Data_43 <= verilogPut_Data_3_21;
              end
            endcase
          end
          else begin
            verilogPut_Found_40 <= 0;
            case (verilogPut_size_3)
              0: begin
                verilogPut_StuckIndex_45 <= 0;
                verilogPut_Data_43 <= verilogPut_Data_0_9;
              end
              1: begin
                verilogPut_StuckIndex_45 <= 1;
                verilogPut_Data_43 <= verilogPut_Data_1_13;
              end
              2: begin
                verilogPut_StuckIndex_45 <= 2;
                verilogPut_Data_43 <= verilogPut_Data_2_17;
              end
              3: begin
                verilogPut_StuckIndex_45 <= 3;
                verilogPut_Data_43 <= verilogPut_Data_3_21;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        209: begin
          verilogPut_child_101 <= verilogPut_Data_43;
          verilogPut_childInparent_103 <= verilogPut_StuckIndex_45;
          verilogPut_found_104 <= verilogPut_Found_40;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        210: begin
          verilogPut_index_47 <= verilogPut_child_101;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        211: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_47;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_47;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_47;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_47;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        212: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        213: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        214: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        215: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        216: begin
          verilogPut_size_48 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_49 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_51 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_54 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_55 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_58 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_59 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_62 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_63 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_66 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        217: begin
          if (verilogPut_isLeaf_49 == 0) begin
            verilogPut_pc <= 356;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        218: begin
          verilogPut_full_105 <= verilogPut_size_48>=4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        219: begin
          if (verilogPut_full_105 == 0) begin
            verilogPut_pc <= 315;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        220: begin
          if (verilogPut_found_104 == 0) begin
            verilogPut_pc <= 267;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        221: begin
          verilogPut_index_299 <= verilogPut_parent_102;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        222: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_299;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_299;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_299;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_299;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        223: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        224: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        225: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        226: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        227: begin
          verilogPut_size_300 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_301 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_303 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_306 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_307 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_310 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_311 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_314 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_315 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_318 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        228: begin
          case (verilogPut_childInparent_103)
            0: begin
              verilogPut_childKey_407 <= verilogPut_Key_0_303;
              verilogPut_childData_408 <= verilogPut_Data_0_306;
            end
            1: begin
              verilogPut_childKey_407 <= verilogPut_Key_1_307;
              verilogPut_childData_408 <= verilogPut_Data_1_310;
            end
            2: begin
              verilogPut_childKey_407 <= verilogPut_Key_2_311;
              verilogPut_childData_408 <= verilogPut_Data_2_314;
            end
            3: begin
              verilogPut_childKey_407 <= verilogPut_Key_3_315;
              verilogPut_childData_408 <= verilogPut_Data_3_318;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        229: begin
          verilogPut_index_326 <= verilogPut_childData_408;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        230: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_326;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_326;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_326;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_326;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        231: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        232: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        233: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        234: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        235: begin
          verilogPut_size_327 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_328 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_330 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_333 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_334 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_337 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_338 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_341 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_342 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_345 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        236: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        237: begin
          verilogPut_Key_0_357 <= verilogPut_Key_0_330;
          verilogPut_Data_0_360 <= verilogPut_Data_0_333;
          verilogPut_Key_1_361 <= verilogPut_Key_1_334;
          verilogPut_Data_1_364 <= verilogPut_Data_1_337;
          verilogPut_size_354 <= 2;
          verilogPut_Key_0_330 <= verilogPut_Key_2_338;
          verilogPut_Data_0_333 <= verilogPut_Data_2_341;
          verilogPut_Key_1_334 <= verilogPut_Key_3_342;
          verilogPut_Data_1_337 <= verilogPut_Data_3_345;
          verilogPut_size_327 <= 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        238: begin
          verilogPut_root_412 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        239: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_412;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        240: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        241: begin
          verilogPut_indexLeft_409 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        242: begin
          if (verilogPut_indexLeft_409 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_414 <= 1;
          verilogPut_isFree_415 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        243: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexLeft_409;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexLeft_409;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_414;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_409;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_415;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        244: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        245: begin
          verilogPut_next_413 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        246: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_412;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_413;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        247: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        248: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        249: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        250: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_childData_408;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_327;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_childData_408;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_330;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_334;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_338;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_342;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_childData_408;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_333;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_337;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_341;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_345;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        251: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        252: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        253: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        254: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexLeft_409;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_354;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexLeft_409;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_357;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_361;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_365;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_369;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexLeft_409;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_360;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_364;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_368;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_372;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        255: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        256: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        257: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        258: begin
          case (verilogPut_size_354)
            1: begin
              verilogPut_Key_374 <= verilogPut_Key_0_357;
              verilogPut_Data_376 <= verilogPut_Data_0_360;
            end
            2: begin
              verilogPut_Key_374 <= verilogPut_Key_1_361;
              verilogPut_Data_376 <= verilogPut_Data_1_364;
            end
            3: begin
              verilogPut_Key_374 <= verilogPut_Key_2_365;
              verilogPut_Data_376 <= verilogPut_Data_2_368;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        259: begin
          verilogPut_Key_347 <= verilogPut_Key_0_330;
          verilogPut_Data_349 <= verilogPut_Data_0_333;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        260: begin
          verilogPut_midKey_411 <= (verilogPut_Key_374 + verilogPut_Key_347) / 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        261: begin
          verilogPut_size_300 <= verilogPut_size_300+1;
          if (3 > verilogPut_childInparent_103) begin
            verilogPut_Key_3_315 <= verilogPut_Key_2_311;
            verilogPut_Data_3_318 <= verilogPut_Data_2_314;
          end
          if (2 > verilogPut_childInparent_103) begin
            verilogPut_Key_2_311 <= verilogPut_Key_1_307;
            verilogPut_Data_2_314 <= verilogPut_Data_1_310;
          end
          if (1 > verilogPut_childInparent_103) begin
            verilogPut_Key_1_307 <= verilogPut_Key_0_303;
            verilogPut_Data_1_310 <= verilogPut_Data_0_306;
          end
          case (verilogPut_childInparent_103)
            0: begin
              verilogPut_Key_0_303 <= verilogPut_midKey_411;
              verilogPut_Data_0_306 <= verilogPut_indexLeft_409;
            end
            1: begin
              verilogPut_Key_1_307 <= verilogPut_midKey_411;
              verilogPut_Data_1_310 <= verilogPut_indexLeft_409;
            end
            2: begin
              verilogPut_Key_2_311 <= verilogPut_midKey_411;
              verilogPut_Data_2_314 <= verilogPut_indexLeft_409;
            end
            3: begin
              verilogPut_Key_3_315 <= verilogPut_midKey_411;
              verilogPut_Data_3_318 <= verilogPut_indexLeft_409;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        262: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_299;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_300;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_299;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_303;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_307;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_311;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_315;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_299;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_306;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_310;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_314;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_318;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        263: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        264: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        265: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        266: begin
          verilogPut_pc <= 314;
        end
        267: begin
          verilogPut_index_416 <= verilogPut_parent_102;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        268: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_416;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_416;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_416;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_416;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        269: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        270: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        271: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        272: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        273: begin
          verilogPut_size_417 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_418 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_420 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_423 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_424 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_427 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_428 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_431 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_432 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_435 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        274: begin
          case (verilogPut_size_417)
            0: begin
              verilogPut_Key_437 <= verilogPut_Key_0_420;
              verilogPut_Data_439 <= verilogPut_Data_0_423;
            end
            1: begin
              verilogPut_Key_437 <= verilogPut_Key_1_424;
              verilogPut_Data_439 <= verilogPut_Data_1_427;
            end
            2: begin
              verilogPut_Key_437 <= verilogPut_Key_2_428;
              verilogPut_Data_439 <= verilogPut_Data_2_431;
            end
            3: begin
              verilogPut_Key_437 <= verilogPut_Key_3_432;
              verilogPut_Data_439 <= verilogPut_Data_3_435;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        275: begin
          verilogPut_childIndex_497 <= verilogPut_Data_439;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        276: begin
          verilogPut_index_443 <= verilogPut_childIndex_497;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        277: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_443;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_443;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_443;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_443;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        278: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        279: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        280: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        281: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        282: begin
          verilogPut_size_444 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_445 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_447 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_450 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_451 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_454 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_455 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_458 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_459 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_462 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        283: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        284: begin
          verilogPut_Key_0_474 <= verilogPut_Key_0_447;
          verilogPut_Data_0_477 <= verilogPut_Data_0_450;
          verilogPut_Key_1_478 <= verilogPut_Key_1_451;
          verilogPut_Data_1_481 <= verilogPut_Data_1_454;
          verilogPut_size_471 <= 2;
          verilogPut_Key_0_447 <= verilogPut_Key_2_455;
          verilogPut_Data_0_450 <= verilogPut_Data_2_458;
          verilogPut_Key_1_451 <= verilogPut_Key_3_459;
          verilogPut_Data_1_454 <= verilogPut_Data_3_462;
          verilogPut_size_444 <= 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        285: begin
          verilogPut_root_500 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        286: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_500;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        287: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        288: begin
          verilogPut_leftIndex_498 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        289: begin
          if (verilogPut_leftIndex_498 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_502 <= 1;
          verilogPut_isFree_503 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        290: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_leftIndex_498;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_leftIndex_498;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_502;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_leftIndex_498;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_503;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        291: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        292: begin
          verilogPut_next_501 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        293: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_500;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_501;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        294: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        295: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        296: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        297: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_leftIndex_498;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_471;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_leftIndex_498;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_474;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_478;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_482;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_486;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_leftIndex_498;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_477;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_481;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_485;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_489;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        298: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        299: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        300: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        301: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_childIndex_497;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_444;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_childIndex_497;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_447;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_451;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_455;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_459;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_childIndex_497;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_450;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_454;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_458;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_462;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        302: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        303: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        304: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        305: begin
          case (verilogPut_size_471)
            1: begin
              verilogPut_Key_491 <= verilogPut_Key_0_474;
              verilogPut_Data_493 <= verilogPut_Data_0_477;
            end
            2: begin
              verilogPut_Key_491 <= verilogPut_Key_1_478;
              verilogPut_Data_493 <= verilogPut_Data_1_481;
            end
            3: begin
              verilogPut_Key_491 <= verilogPut_Key_2_482;
              verilogPut_Data_493 <= verilogPut_Data_2_485;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        306: begin
          verilogPut_Key_464 <= verilogPut_Key_0_447;
          verilogPut_Data_466 <= verilogPut_Data_0_450;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        307: begin
          verilogPut_midKey_499 <= (verilogPut_Key_491 + verilogPut_Key_464) / 2;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        308: begin
          case (verilogPut_size_417)
            0: begin
              verilogPut_Key_0_420 <= verilogPut_midKey_499;
              verilogPut_Data_0_423 <= verilogPut_leftIndex_498;
            end
            1: begin
              verilogPut_Key_1_424 <= verilogPut_midKey_499;
              verilogPut_Data_1_427 <= verilogPut_leftIndex_498;
            end
            2: begin
              verilogPut_Key_2_428 <= verilogPut_midKey_499;
              verilogPut_Data_2_431 <= verilogPut_leftIndex_498;
            end
            3: begin
              verilogPut_Key_3_432 <= verilogPut_midKey_499;
              verilogPut_Data_3_435 <= verilogPut_leftIndex_498;
            end
          endcase
          verilogPut_size_417 <= verilogPut_size_417+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        309: begin
          case (verilogPut_size_417)
            0: begin
              verilogPut_Key_0_420 <= verilogPut_midKey_499;
              verilogPut_Data_0_423 <= verilogPut_childIndex_497;
            end
            1: begin
              verilogPut_Key_1_424 <= verilogPut_midKey_499;
              verilogPut_Data_1_427 <= verilogPut_childIndex_497;
            end
            2: begin
              verilogPut_Key_2_428 <= verilogPut_midKey_499;
              verilogPut_Data_2_431 <= verilogPut_childIndex_497;
            end
            3: begin
              verilogPut_Key_3_432 <= verilogPut_midKey_499;
              verilogPut_Data_3_435 <= verilogPut_childIndex_497;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        310: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_416;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_417;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_416;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_420;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_424;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_428;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_432;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_416;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_423;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_427;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_431;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_435;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        311: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        312: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        313: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        314: begin
          verilogPut_pc <= 315;
        end
        315: begin
          verilogPut_BtreeIndex_98 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        316: begin
          verilogPut_index_74 <= verilogPut_BtreeIndex_98;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        317: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_74;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_74;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_74;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_74;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        318: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        319: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        320: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        321: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        322: begin
          verilogPut_size_75 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_76 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_78 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_81 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_82 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_85 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_86 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_89 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_90 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_93 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        323: begin
          if (verilogPut_isLeaf_76 == 0) begin
            verilogPut_pc <= 330;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        324: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 == verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 == verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 == verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 == verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        325: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        326: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        327: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Key_95 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Key_95 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Key_95 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Key_95 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        328: begin
          verilogPut_pc <= 336;
        end
        329: begin
          verilogPut_pc <= 336;
        end
        330: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 <= verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 >  verilogPut_Key_0_78 && verilogPut_k_0 <= verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 >  verilogPut_Key_1_82 && verilogPut_k_0 <= verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 >  verilogPut_Key_2_86 && verilogPut_k_0 <= verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        331: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        332: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        333: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_FoundKey_96 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_FoundKey_96 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_FoundKey_96 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_FoundKey_96 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
            case (verilogPut_size_75)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        334: begin
          verilogPut_BtreeIndex_98 <= verilogPut_Data_97;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        335: begin
          verilogPut_pc <= 316;
        end
        336: begin
          if (verilogPut_Found_94 == 0) begin
            verilogPut_pc <= 339;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        337: begin
          if (verilogPut_StuckIndex_99 == verilogPut_size_75) begin
            verilogPut_size_75 <= verilogPut_size_75+1;
          end
          case (verilogPut_StuckIndex_99)
            0: begin
              verilogPut_Key_0_78 <= verilogPut_k_0;
              verilogPut_Data_0_81 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_82 <= verilogPut_k_0;
              verilogPut_Data_1_85 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_86 <= verilogPut_k_0;
              verilogPut_Data_2_89 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_90 <= verilogPut_k_0;
              verilogPut_Data_3_93 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        338: begin
          verilogPut_pc <= 350;
        end
        339: begin
          verilogPut_notFull_505 <= verilogPut_size_75< 4 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        340: begin
          if (verilogPut_notFull_505 == 0) begin
            verilogPut_pc <= 349;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        341: begin
          verilogPut_KeyCompares_0_79 <= verilogPut_k_0 <= verilogPut_Key_0_78 && 0 < verilogPut_size_75;
          verilogPut_KeyCollapse_0_80 <= 0;
          verilogPut_KeyCompares_1_83 <= verilogPut_k_0 >  verilogPut_Key_0_78 && verilogPut_k_0 <= verilogPut_Key_1_82 && 1 < verilogPut_size_75;
          verilogPut_KeyCollapse_1_84 <= 1;
          verilogPut_KeyCompares_2_87 <= verilogPut_k_0 >  verilogPut_Key_1_82 && verilogPut_k_0 <= verilogPut_Key_2_86 && 2 < verilogPut_size_75;
          verilogPut_KeyCollapse_2_88 <= 2;
          verilogPut_KeyCompares_3_91 <= verilogPut_k_0 >  verilogPut_Key_2_86 && verilogPut_k_0 <= verilogPut_Key_3_90 && 3 < verilogPut_size_75;
          verilogPut_KeyCollapse_3_92 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        342: begin
          if (verilogPut_KeyCompares_1_83) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_1_84;
          end
          if (verilogPut_KeyCompares_3_91) begin
            verilogPut_KeyCompares_2_87 <= 1;
            verilogPut_KeyCollapse_2_88 <= verilogPut_KeyCollapse_3_92;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        343: begin
          if (verilogPut_KeyCompares_2_87) begin
            verilogPut_KeyCompares_0_79 <= 1;
            verilogPut_KeyCollapse_0_80 <= verilogPut_KeyCollapse_2_88;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        344: begin
          if (verilogPut_KeyCompares_0_79) begin
            verilogPut_Found_94 <= 1;
            case (verilogPut_KeyCollapse_0_80)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_FoundKey_96 <= verilogPut_Key_0_78;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_FoundKey_96 <= verilogPut_Key_1_82;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_FoundKey_96 <= verilogPut_Key_2_86;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_FoundKey_96 <= verilogPut_Key_3_90;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          else begin
            verilogPut_Found_94 <= 0;
            case (verilogPut_size_75)
              0: begin
                verilogPut_StuckIndex_99 <= 0;
                verilogPut_Data_97 <= verilogPut_Data_0_81;
              end
              1: begin
                verilogPut_StuckIndex_99 <= 1;
                verilogPut_Data_97 <= verilogPut_Data_1_85;
              end
              2: begin
                verilogPut_StuckIndex_99 <= 2;
                verilogPut_Data_97 <= verilogPut_Data_2_89;
              end
              3: begin
                verilogPut_StuckIndex_99 <= 3;
                verilogPut_Data_97 <= verilogPut_Data_3_93;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        345: begin
          verilogPut_size_75 <= verilogPut_size_75+1;
          if (3 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_3_90 <= verilogPut_Key_2_86;
            verilogPut_Data_3_93 <= verilogPut_Data_2_89;
          end
          if (2 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_2_86 <= verilogPut_Key_1_82;
            verilogPut_Data_2_89 <= verilogPut_Data_1_85;
          end
          if (1 > verilogPut_StuckIndex_99) begin
            verilogPut_Key_1_82 <= verilogPut_Key_0_78;
            verilogPut_Data_1_85 <= verilogPut_Data_0_81;
          end
          case (verilogPut_StuckIndex_99)
            0: begin
              verilogPut_Key_0_78 <= verilogPut_k_0;
              verilogPut_Data_0_81 <= verilogPut_d_1;
            end
            1: begin
              verilogPut_Key_1_82 <= verilogPut_k_0;
              verilogPut_Data_1_85 <= verilogPut_d_1;
            end
            2: begin
              verilogPut_Key_2_86 <= verilogPut_k_0;
              verilogPut_Data_2_89 <= verilogPut_d_1;
            end
            3: begin
              verilogPut_Key_3_90 <= verilogPut_k_0;
              verilogPut_Data_3_93 <= verilogPut_d_1;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        346: begin
          verilogPut_Found_94 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        347: begin
          verilogPut_pc <= verilogPut_pc + 1;
        end
        348: begin
          verilogPut_pc <= 350;
        end
        349: begin
          verilogPut_pc <= 354;
        end
        350: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_74;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_75;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_74;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_78;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_82;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_86;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_90;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_74;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_81;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_85;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_89;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_93;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        351: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        352: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        353: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        354: begin
          verilogPut_pc <= 449;
        end
        355: begin
          verilogPut_pc <= 449;
        end
        356: begin
          verilogPut_full_105 <= verilogPut_size_48>=3 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        357: begin
          if (verilogPut_full_105 == 0) begin
            verilogPut_pc <= 447;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        358: begin
          if (verilogPut_found_104 == 0) begin
            verilogPut_pc <= 402;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        359: begin
          verilogPut_index_506 <= verilogPut_parent_102;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        360: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_506;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_506;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_506;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_506;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        361: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        362: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        363: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        364: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        365: begin
          verilogPut_size_507 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_508 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_510 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_513 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_514 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_517 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_518 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_521 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_522 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_525 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        366: begin
          case (verilogPut_childInparent_103)
            0: begin
              verilogPut_childKey_614 <= verilogPut_Key_0_510;
              verilogPut_childData_615 <= verilogPut_Data_0_513;
            end
            1: begin
              verilogPut_childKey_614 <= verilogPut_Key_1_514;
              verilogPut_childData_615 <= verilogPut_Data_1_517;
            end
            2: begin
              verilogPut_childKey_614 <= verilogPut_Key_2_518;
              verilogPut_childData_615 <= verilogPut_Data_2_521;
            end
            3: begin
              verilogPut_childKey_614 <= verilogPut_Key_3_522;
              verilogPut_childData_615 <= verilogPut_Data_3_525;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        367: begin
          verilogPut_index_533 <= verilogPut_childData_615;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        368: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_533;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_533;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_533;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_533;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        369: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        370: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        371: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        372: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        373: begin
          verilogPut_size_534 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_535 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_537 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_540 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_541 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_544 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_545 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_548 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_549 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_552 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        374: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        375: begin
          verilogPut_Key_0_564 <= verilogPut_Key_0_537;
          verilogPut_Data_0_567 <= verilogPut_Data_0_540;
          verilogPut_size_561 <= 1;
          verilogPut_Data_1_571 <= verilogPut_Data_1_544;
          verilogPut_childKey_614 <= verilogPut_Key_1_541;
          verilogPut_Key_0_537 <= verilogPut_Key_2_545;
          verilogPut_Data_0_540 <= verilogPut_Data_2_548;
          verilogPut_Key_1_541 <= verilogPut_Key_3_549;
          verilogPut_Data_1_544 <= verilogPut_Data_3_552;
          verilogPut_size_534 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        376: begin
          verilogPut_root_619 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        377: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_619;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        378: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        379: begin
          verilogPut_indexLeft_616 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        380: begin
          if (verilogPut_indexLeft_616 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_621 <= 0;
          verilogPut_isFree_622 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        381: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexLeft_616;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexLeft_616;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_621;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_616;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_622;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        382: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        383: begin
          verilogPut_next_620 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        384: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_619;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_620;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        385: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        386: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        387: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        388: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexLeft_616;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_561;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexLeft_616;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_564;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_568;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_572;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_576;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexLeft_616;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_567;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_571;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_575;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_579;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        389: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        390: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        391: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        392: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_childData_615;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_534;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_childData_615;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_537;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_541;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_545;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_549;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_childData_615;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_540;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_544;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_548;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_552;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        393: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        394: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        395: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        396: begin
          verilogPut_size_507 <= verilogPut_size_507+1;
          if (3 > verilogPut_childInparent_103) begin
            verilogPut_Key_3_522 <= verilogPut_Key_2_518;
            verilogPut_Data_3_525 <= verilogPut_Data_2_521;
          end
          if (2 > verilogPut_childInparent_103) begin
            verilogPut_Key_2_518 <= verilogPut_Key_1_514;
            verilogPut_Data_2_521 <= verilogPut_Data_1_517;
          end
          if (1 > verilogPut_childInparent_103) begin
            verilogPut_Key_1_514 <= verilogPut_Key_0_510;
            verilogPut_Data_1_517 <= verilogPut_Data_0_513;
          end
          case (verilogPut_childInparent_103)
            0: begin
              verilogPut_Key_0_510 <= verilogPut_childKey_614;
              verilogPut_Data_0_513 <= verilogPut_indexLeft_616;
            end
            1: begin
              verilogPut_Key_1_514 <= verilogPut_childKey_614;
              verilogPut_Data_1_517 <= verilogPut_indexLeft_616;
            end
            2: begin
              verilogPut_Key_2_518 <= verilogPut_childKey_614;
              verilogPut_Data_2_521 <= verilogPut_indexLeft_616;
            end
            3: begin
              verilogPut_Key_3_522 <= verilogPut_childKey_614;
              verilogPut_Data_3_525 <= verilogPut_indexLeft_616;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        397: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_506;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_507;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_506;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_510;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_514;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_518;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_522;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_506;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_513;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_517;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_521;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_525;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        398: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        399: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        400: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        401: begin
          verilogPut_pc <= 446;
        end
        402: begin
          verilogPut_index_623 <= verilogPut_parent_102;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        403: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_623;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_623;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_623;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_623;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        404: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        405: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        406: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        407: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        408: begin
          verilogPut_size_624 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_625 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_627 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_630 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_631 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_634 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_635 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_638 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_639 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_642 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        409: begin
          case (verilogPut_size_624)
            0: begin
              verilogPut_Key_644 <= verilogPut_Key_0_627;
              verilogPut_Data_646 <= verilogPut_Data_0_630;
            end
            1: begin
              verilogPut_Key_644 <= verilogPut_Key_1_631;
              verilogPut_Data_646 <= verilogPut_Data_1_634;
            end
            2: begin
              verilogPut_Key_644 <= verilogPut_Key_2_635;
              verilogPut_Data_646 <= verilogPut_Data_2_638;
            end
            3: begin
              verilogPut_Key_644 <= verilogPut_Key_3_639;
              verilogPut_Data_646 <= verilogPut_Data_3_642;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        410: begin
          verilogPut_childData_732 <= verilogPut_Data_646;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        411: begin
          verilogPut_index_650 <= verilogPut_childData_732;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        412: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_650;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_650;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_650;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_650;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        413: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        414: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        415: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        416: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        417: begin
          verilogPut_size_651 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_652 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_654 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_657 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_658 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_661 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_662 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_665 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_666 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_669 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        418: begin
          
          verilogPut_pc <= verilogPut_pc + 1;
        end
        419: begin
          verilogPut_Key_0_681 <= verilogPut_Key_0_654;
          verilogPut_Data_0_684 <= verilogPut_Data_0_657;
          verilogPut_size_678 <= 1;
          verilogPut_Data_1_688 <= verilogPut_Data_1_661;
          verilogPut_midKey_735 <= verilogPut_Key_1_658;
          verilogPut_Key_0_654 <= verilogPut_Key_2_662;
          verilogPut_Data_0_657 <= verilogPut_Data_2_665;
          verilogPut_Key_1_658 <= verilogPut_Key_3_666;
          verilogPut_Data_1_661 <= verilogPut_Data_3_669;
          verilogPut_size_651 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        420: begin
          verilogPut_root_736 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        421: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_736;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        422: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        423: begin
          verilogPut_indexLeft_733 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        424: begin
          if (verilogPut_indexLeft_733 == 0) begin
            verilogPut_returnCode <= 20;
            verilogPut_stop <= 1;
          end
          verilogPut_isLeaf_738 <= 0;
          verilogPut_isFree_739 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        425: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_indexLeft_733;
          freeNext_9_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_indexLeft_733;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_738;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_733;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_739;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        426: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        427: begin
          verilogPut_next_737 <= freeNext_freeNext_9_result_0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        428: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_root_736;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_737;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        429: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        430: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        431: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        432: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_indexLeft_733;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_678;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_indexLeft_733;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_681;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_685;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_689;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_693;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_indexLeft_733;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_684;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_688;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_692;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_696;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        433: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        434: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        435: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        436: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_childData_732;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_651;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_childData_732;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_654;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_658;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_662;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_666;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_childData_732;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_657;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_661;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_665;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_669;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        437: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        438: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        439: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        440: begin
          case (verilogPut_size_624)
            0: begin
              verilogPut_Key_0_627 <= verilogPut_midKey_735;
              verilogPut_Data_0_630 <= verilogPut_indexLeft_733;
            end
            1: begin
              verilogPut_Key_1_631 <= verilogPut_midKey_735;
              verilogPut_Data_1_634 <= verilogPut_indexLeft_733;
            end
            2: begin
              verilogPut_Key_2_635 <= verilogPut_midKey_735;
              verilogPut_Data_2_638 <= verilogPut_indexLeft_733;
            end
            3: begin
              verilogPut_Key_3_639 <= verilogPut_midKey_735;
              verilogPut_Data_3_642 <= verilogPut_indexLeft_733;
            end
          endcase
          verilogPut_size_624 <= verilogPut_size_624+1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        441: begin
          case (verilogPut_size_624)
            0: begin
              verilogPut_Key_0_627 <= verilogPut_midKey_735;
              verilogPut_Data_0_630 <= verilogPut_childData_732;
            end
            1: begin
              verilogPut_Key_1_631 <= verilogPut_midKey_735;
              verilogPut_Data_1_634 <= verilogPut_childData_732;
            end
            2: begin
              verilogPut_Key_2_635 <= verilogPut_midKey_735;
              verilogPut_Data_2_638 <= verilogPut_childData_732;
            end
            3: begin
              verilogPut_Key_3_639 <= verilogPut_midKey_735;
              verilogPut_Data_3_642 <= verilogPut_childData_732;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        442: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_623;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_624;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_623;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_627;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_631;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_635;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_639;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_623;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_630;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_634;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_638;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_642;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        443: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        444: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        445: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        446: begin
          verilogPut_pc <= 448;
        end
        447: begin
          verilogPut_parent_102 <= verilogPut_child_101;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        448: begin
          verilogPut_pc <= 198;
        end
        449: begin
          verilogPut_position_767 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        450: begin
          verilogPut_index_740 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        451: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        452: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        453: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        454: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        455: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        456: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        457: begin
          if (verilogPut_isLeaf_742 == 0) begin
            verilogPut_pc <= 460;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        458: begin
          verilogPut_pc <= 1000;
        end
        459: begin
          verilogPut_pc <= 460;
        end
        460: begin
          verilogPut_success_857 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        461: begin
          verilogPut_index_771 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        462: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_771;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_771;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_771;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_771;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        463: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        464: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        465: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        466: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        467: begin
          verilogPut_size_772 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_773 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_775 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_778 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_779 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_782 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_783 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_786 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_787 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_790 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        468: begin
          verilogPut_test_858 <= verilogPut_size_772==1 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        469: begin
          if (verilogPut_test_858 == 0) begin
            verilogPut_pc <= 521;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        470: begin
          verilogPut_indexLeft_854 <= verilogPut_Data_0_778;
          verilogPut_indexRight_855 <= verilogPut_Data_1_782;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        471: begin
          verilogPut_index_798 <= verilogPut_indexLeft_854;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        472: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_798;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_798;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_798;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_798;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        473: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        474: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        475: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        476: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        477: begin
          verilogPut_size_799 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_800 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_802 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_805 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_806 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_809 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_810 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_813 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_814 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_817 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        478: begin
          verilogPut_index_825 <= verilogPut_indexRight_855;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        479: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_825;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_825;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_825;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_825;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        480: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        481: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        482: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        483: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        484: begin
          verilogPut_size_826 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_827 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_829 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_832 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_833 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_836 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_837 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_840 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_841 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_844 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        485: begin
          if (verilogPut_isLeaf_800 == 0) begin
            verilogPut_pc <= 521;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        486: begin
          if (verilogPut_isLeaf_827 == 0) begin
            verilogPut_pc <= 520;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        487: begin
          verilogPut_MergeSuccess_797 <= 0;
          case (verilogPut_size_799)
            0: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                4: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        488: begin
          if (verilogPut_MergeSuccess_797 == 0) begin
            verilogPut_pc <= 492;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        489: begin
          verilogPut_MergeSuccess_797 <= 0;
          case (verilogPut_size_772)
            0: begin
              case (verilogPut_size_799)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_802;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_805;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_802;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_805;
                  verilogPut_Key_1_779 <= verilogPut_Key_1_806;
                  verilogPut_Data_1_782 <= verilogPut_Data_1_809;
                  verilogPut_size_772 <= verilogPut_size_772 + 2;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_802;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_805;
                  verilogPut_Key_1_779 <= verilogPut_Key_1_806;
                  verilogPut_Data_1_782 <= verilogPut_Data_1_809;
                  verilogPut_Key_2_783 <= verilogPut_Key_2_810;
                  verilogPut_Data_2_786 <= verilogPut_Data_2_813;
                  verilogPut_size_772 <= verilogPut_size_772 + 3;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                4: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_802;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_805;
                  verilogPut_Key_1_779 <= verilogPut_Key_1_806;
                  verilogPut_Data_1_782 <= verilogPut_Data_1_809;
                  verilogPut_Key_2_783 <= verilogPut_Key_2_810;
                  verilogPut_Data_2_786 <= verilogPut_Data_2_813;
                  verilogPut_Key_3_787 <= verilogPut_Key_3_814;
                  verilogPut_Data_3_790 <= verilogPut_Data_3_817;
                  verilogPut_size_772 <= verilogPut_size_772 + 4;
                  verilogPut_MergeSuccess_797 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_799)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_1_779 <= verilogPut_Key_0_802;
                  verilogPut_Data_1_782 <= verilogPut_Data_0_805;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_Key_1_779 <= verilogPut_Key_0_802;
                  verilogPut_Data_1_782 <= verilogPut_Data_0_805;
                  verilogPut_Key_2_783 <= verilogPut_Key_1_806;
                  verilogPut_Data_2_786 <= verilogPut_Data_1_809;
                  verilogPut_size_772 <= verilogPut_size_772 + 2;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                  verilogPut_Key_1_779 <= verilogPut_Key_0_802;
                  verilogPut_Data_1_782 <= verilogPut_Data_0_805;
                  verilogPut_Key_2_783 <= verilogPut_Key_1_806;
                  verilogPut_Data_2_786 <= verilogPut_Data_1_809;
                  verilogPut_Key_3_787 <= verilogPut_Key_2_810;
                  verilogPut_Data_3_790 <= verilogPut_Data_2_813;
                  verilogPut_size_772 <= verilogPut_size_772 + 3;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_799)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_2_783 <= verilogPut_Key_0_802;
                  verilogPut_Data_2_786 <= verilogPut_Data_0_805;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_Key_2_783 <= verilogPut_Key_0_802;
                  verilogPut_Data_2_786 <= verilogPut_Data_0_805;
                  verilogPut_Key_3_787 <= verilogPut_Key_1_806;
                  verilogPut_Data_3_790 <= verilogPut_Data_1_809;
                  verilogPut_size_772 <= verilogPut_size_772 + 2;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_799)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_3_787 <= verilogPut_Key_0_802;
                  verilogPut_Data_3_790 <= verilogPut_Data_0_805;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_799)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        490: begin
          verilogPut_MergeSuccess_797 <= 0;
          case (verilogPut_size_772)
            0: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_829;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_832;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_829;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_832;
                  verilogPut_Key_1_779 <= verilogPut_Key_1_833;
                  verilogPut_Data_1_782 <= verilogPut_Data_1_836;
                  verilogPut_size_772 <= verilogPut_size_772 + 2;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_829;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_832;
                  verilogPut_Key_1_779 <= verilogPut_Key_1_833;
                  verilogPut_Data_1_782 <= verilogPut_Data_1_836;
                  verilogPut_Key_2_783 <= verilogPut_Key_2_837;
                  verilogPut_Data_2_786 <= verilogPut_Data_2_840;
                  verilogPut_size_772 <= verilogPut_size_772 + 3;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                4: begin
                  verilogPut_Key_0_775 <= verilogPut_Key_0_829;
                  verilogPut_Data_0_778 <= verilogPut_Data_0_832;
                  verilogPut_Key_1_779 <= verilogPut_Key_1_833;
                  verilogPut_Data_1_782 <= verilogPut_Data_1_836;
                  verilogPut_Key_2_783 <= verilogPut_Key_2_837;
                  verilogPut_Data_2_786 <= verilogPut_Data_2_840;
                  verilogPut_Key_3_787 <= verilogPut_Key_3_841;
                  verilogPut_Data_3_790 <= verilogPut_Data_3_844;
                  verilogPut_size_772 <= verilogPut_size_772 + 4;
                  verilogPut_MergeSuccess_797 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_1_779 <= verilogPut_Key_0_829;
                  verilogPut_Data_1_782 <= verilogPut_Data_0_832;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_Key_1_779 <= verilogPut_Key_0_829;
                  verilogPut_Data_1_782 <= verilogPut_Data_0_832;
                  verilogPut_Key_2_783 <= verilogPut_Key_1_833;
                  verilogPut_Data_2_786 <= verilogPut_Data_1_836;
                  verilogPut_size_772 <= verilogPut_size_772 + 2;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                  verilogPut_Key_1_779 <= verilogPut_Key_0_829;
                  verilogPut_Data_1_782 <= verilogPut_Data_0_832;
                  verilogPut_Key_2_783 <= verilogPut_Key_1_833;
                  verilogPut_Data_2_786 <= verilogPut_Data_1_836;
                  verilogPut_Key_3_787 <= verilogPut_Key_2_837;
                  verilogPut_Data_3_790 <= verilogPut_Data_2_840;
                  verilogPut_size_772 <= verilogPut_size_772 + 3;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_2_783 <= verilogPut_Key_0_829;
                  verilogPut_Data_2_786 <= verilogPut_Data_0_832;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                  verilogPut_Key_2_783 <= verilogPut_Key_0_829;
                  verilogPut_Data_2_786 <= verilogPut_Data_0_832;
                  verilogPut_Key_3_787 <= verilogPut_Key_1_833;
                  verilogPut_Data_3_790 <= verilogPut_Data_1_836;
                  verilogPut_size_772 <= verilogPut_size_772 + 2;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                  verilogPut_Key_3_787 <= verilogPut_Key_0_829;
                  verilogPut_Data_3_790 <= verilogPut_Data_0_832;
                  verilogPut_size_772 <= verilogPut_size_772 + 1;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_826)
                0: begin
                  verilogPut_size_772 <= verilogPut_size_772 + 0;
                  verilogPut_MergeSuccess_797 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        491: begin
          verilogPut_pc <= 492;
        end
        492: begin
          if (verilogPut_MergeSuccess_797 == 0) begin
            verilogPut_pc <= 519;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        493: begin
          verilogPut_isLeaf_773 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        494: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_771;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_772;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckIsLeaf_8_index_38 <= verilogPut_index_771;
          verilogPut_stuckIsLeaf_8_value_39 <= verilogPut_isLeaf_773;
          stuckIsLeaf_8_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_771;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_775;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_779;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_783;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_787;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_771;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_778;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_782;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_786;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_790;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        495: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        496: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        497: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        498: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        499: begin
          verilogPut_root_860 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        500: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_860;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        501: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        502: begin
          verilogPut_next_859 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_860;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexLeft_854;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_861 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        503: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_854;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_861;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        504: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        505: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexLeft_854;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_859;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        506: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        507: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        508: begin
          verilogPut_root_863 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        509: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_863;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        510: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        511: begin
          verilogPut_next_862 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_863;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_855;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_864 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        512: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_855;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_864;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        513: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        514: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_855;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_862;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        515: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        516: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        517: begin
          verilogPut_success_857 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        518: begin
          verilogPut_pc <= 519;
        end
        519: begin
          verilogPut_pc <= 520;
        end
        520: begin
          verilogPut_pc <= 521;
        end
        521: begin
          if (verilogPut_success_857 == 0) begin
            verilogPut_pc <= 524;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        522: begin
          verilogPut_pc <= 1000;
        end
        523: begin
          verilogPut_pc <= 524;
        end
        524: begin
          verilogPut_index_865 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        525: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_865;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_865;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_865;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_865;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        526: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        527: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        528: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        529: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        530: begin
          verilogPut_size_866 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_867 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_869 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_872 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_873 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_876 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_877 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_880 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_881 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_884 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        531: begin
          verilogPut_success_953 <= 0;
          if (verilogPut_size_866 != 1) begin
            verilogPut_pc <= 577;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        532: begin
          verilogPut_midKey_952 <= verilogPut_Key_0_869;
          verilogPut_indexLeft_950 <= verilogPut_Data_0_872;
          verilogPut_indexRight_951 <= verilogPut_Data_1_876;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        533: begin
          if (verilogPut_isLeaf_894 == 0) begin
            verilogPut_pc <= 535;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        534: begin
          verilogPut_pc <= 577;
        end
        535: begin
          if (verilogPut_isLeaf_921 == 0) begin
            verilogPut_pc <= 537;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        536: begin
          verilogPut_pc <= 577;
        end
        537: begin
          verilogPut_index_892 <= verilogPut_indexLeft_950;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        538: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_892;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_892;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_892;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_892;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        539: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        540: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        541: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        542: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        543: begin
          verilogPut_size_893 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_894 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_896 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_899 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_900 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_903 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_904 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_907 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_908 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_911 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        544: begin
          verilogPut_index_919 <= verilogPut_indexRight_951;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        545: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_919;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_919;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_919;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_919;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        546: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        547: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        548: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        549: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        550: begin
          verilogPut_size_920 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_921 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_923 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_926 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_927 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_930 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_931 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_934 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_935 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_938 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        551: begin
          verilogPut_MergeSuccess_891 <= 0;
          case (verilogPut_size_893)
            0: begin
              case (verilogPut_size_920)
                0: begin
                  verilogPut_Key_0_869 <= verilogPut_midKey_952;
                  verilogPut_Data_0_872 <= verilogPut_Data_0_899;
                  verilogPut_Data_1_876 <= verilogPut_Data_0_926;
                  verilogPut_size_866 <= 1;
                  verilogPut_MergeSuccess_891 <= 1;
                end
                1: begin
                  verilogPut_Key_0_869 <= verilogPut_midKey_952;
                  verilogPut_Data_0_872 <= verilogPut_Data_0_899;
                  verilogPut_Key_1_873 <= verilogPut_Key_0_923;
                  verilogPut_Data_1_876 <= verilogPut_Data_0_926;
                  verilogPut_Data_2_880 <= verilogPut_Data_1_930;
                  verilogPut_size_866 <= 2;
                  verilogPut_MergeSuccess_891 <= 1;
                end
                2: begin
                  verilogPut_Key_0_869 <= verilogPut_midKey_952;
                  verilogPut_Data_0_872 <= verilogPut_Data_0_899;
                  verilogPut_Key_1_873 <= verilogPut_Key_0_923;
                  verilogPut_Data_1_876 <= verilogPut_Data_0_926;
                  verilogPut_Key_2_877 <= verilogPut_Key_1_927;
                  verilogPut_Data_2_880 <= verilogPut_Data_1_930;
                  verilogPut_Data_3_884 <= verilogPut_Data_2_934;
                  verilogPut_size_866 <= 3;
                  verilogPut_MergeSuccess_891 <= 1;
                end
                3: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_920)
                0: begin
                  verilogPut_Key_0_869 <= verilogPut_Key_0_896;
                  verilogPut_Data_0_872 <= verilogPut_Data_0_899;
                  verilogPut_Key_1_873 <= verilogPut_midKey_952;
                  verilogPut_Data_1_876 <= verilogPut_Data_1_903;
                  verilogPut_Data_2_880 <= verilogPut_Data_0_926;
                  verilogPut_size_866 <= 2;
                  verilogPut_MergeSuccess_891 <= 1;
                end
                1: begin
                  verilogPut_Key_0_869 <= verilogPut_Key_0_896;
                  verilogPut_Data_0_872 <= verilogPut_Data_0_899;
                  verilogPut_Key_1_873 <= verilogPut_midKey_952;
                  verilogPut_Data_1_876 <= verilogPut_Data_1_903;
                  verilogPut_Key_2_877 <= verilogPut_Key_0_923;
                  verilogPut_Data_2_880 <= verilogPut_Data_0_926;
                  verilogPut_Data_3_884 <= verilogPut_Data_1_930;
                  verilogPut_size_866 <= 3;
                  verilogPut_MergeSuccess_891 <= 1;
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_920)
                0: begin
                  verilogPut_Key_0_869 <= verilogPut_Key_0_896;
                  verilogPut_Data_0_872 <= verilogPut_Data_0_899;
                  verilogPut_Key_1_873 <= verilogPut_Key_1_900;
                  verilogPut_Data_1_876 <= verilogPut_Data_1_903;
                  verilogPut_Key_2_877 <= verilogPut_midKey_952;
                  verilogPut_Data_2_880 <= verilogPut_Data_2_907;
                  verilogPut_Data_3_884 <= verilogPut_Data_0_926;
                  verilogPut_size_866 <= 3;
                  verilogPut_MergeSuccess_891 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_920)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        552: begin
          if (verilogPut_MergeSuccess_891 == 0) begin
            verilogPut_pc <= 577;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        553: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_865;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_866;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_865;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_869;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_873;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_877;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_881;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_865;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_872;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_876;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_880;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_884;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        554: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        555: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        556: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        557: begin
          verilogPut_root_956 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        558: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_956;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        559: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        560: begin
          verilogPut_next_955 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_956;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexLeft_950;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_957 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        561: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexLeft_950;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_957;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        562: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        563: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexLeft_950;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_955;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        564: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        565: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        566: begin
          verilogPut_root_959 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        567: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_959;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        568: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        569: begin
          verilogPut_next_958 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_959;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_951;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_960 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        570: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_951;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_960;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        571: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        572: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_951;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_958;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        573: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        574: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        575: begin
          verilogPut_success_953 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        576: begin
          verilogPut_pc <= 577;
        end
        577: begin
          if (verilogPut_success_953 == 0) begin
            verilogPut_pc <= 586;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        578: begin
          verilogPut_index_740 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        579: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        580: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        581: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        582: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        583: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        584: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        585: begin
          verilogPut_pc <= 586;
        end
        586: begin
          verilogPut_success_1021 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        587: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 629;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        588: begin
          verilogPut_size_1016 <= verilogPut_size_741;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        589: begin
          case (verilogPut_size_1016)
            1: begin
              verilogPut_indexLeft_1018 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1019 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_indexLeft_1018 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1019 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_indexLeft_1018 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1019 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        590: begin
          verilogPut_index_961 <= verilogPut_indexLeft_1018;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        591: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_961;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_961;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_961;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_961;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        592: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        593: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        594: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        595: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        596: begin
          verilogPut_size_962 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_963 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_965 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_968 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_969 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_972 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_973 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_976 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_977 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_980 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        597: begin
          verilogPut_index_988 <= verilogPut_indexRight_1019;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        598: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_988;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_988;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_988;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_988;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        599: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        600: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        601: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        602: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        603: begin
          verilogPut_size_989 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_990 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_992 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_995 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_996 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_999 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1000 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1003 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1004 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1007 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        604: begin
          if (verilogPut_isLeaf_963 == 0) begin
            verilogPut_pc <= 629;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        605: begin
          if (verilogPut_isLeaf_990 == 0) begin
            verilogPut_pc <= 628;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        606: begin
          verilogPut_MergeSuccess_987 <= 0;
          case (verilogPut_size_962)
            0: begin
              case (verilogPut_size_989)
                0: begin
                  verilogPut_size_962 <= verilogPut_size_962 + 0;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                1: begin
                  verilogPut_Key_0_965 <= verilogPut_Key_0_992;
                  verilogPut_Data_0_968 <= verilogPut_Data_0_995;
                  verilogPut_size_962 <= verilogPut_size_962 + 1;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                2: begin
                  verilogPut_Key_0_965 <= verilogPut_Key_0_992;
                  verilogPut_Data_0_968 <= verilogPut_Data_0_995;
                  verilogPut_Key_1_969 <= verilogPut_Key_1_996;
                  verilogPut_Data_1_972 <= verilogPut_Data_1_999;
                  verilogPut_size_962 <= verilogPut_size_962 + 2;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                3: begin
                  verilogPut_Key_0_965 <= verilogPut_Key_0_992;
                  verilogPut_Data_0_968 <= verilogPut_Data_0_995;
                  verilogPut_Key_1_969 <= verilogPut_Key_1_996;
                  verilogPut_Data_1_972 <= verilogPut_Data_1_999;
                  verilogPut_Key_2_973 <= verilogPut_Key_2_1000;
                  verilogPut_Data_2_976 <= verilogPut_Data_2_1003;
                  verilogPut_size_962 <= verilogPut_size_962 + 3;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                4: begin
                  verilogPut_Key_0_965 <= verilogPut_Key_0_992;
                  verilogPut_Data_0_968 <= verilogPut_Data_0_995;
                  verilogPut_Key_1_969 <= verilogPut_Key_1_996;
                  verilogPut_Data_1_972 <= verilogPut_Data_1_999;
                  verilogPut_Key_2_973 <= verilogPut_Key_2_1000;
                  verilogPut_Data_2_976 <= verilogPut_Data_2_1003;
                  verilogPut_Key_3_977 <= verilogPut_Key_3_1004;
                  verilogPut_Data_3_980 <= verilogPut_Data_3_1007;
                  verilogPut_size_962 <= verilogPut_size_962 + 4;
                  verilogPut_MergeSuccess_987 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_989)
                0: begin
                  verilogPut_size_962 <= verilogPut_size_962 + 0;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                1: begin
                  verilogPut_Key_1_969 <= verilogPut_Key_0_992;
                  verilogPut_Data_1_972 <= verilogPut_Data_0_995;
                  verilogPut_size_962 <= verilogPut_size_962 + 1;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                2: begin
                  verilogPut_Key_1_969 <= verilogPut_Key_0_992;
                  verilogPut_Data_1_972 <= verilogPut_Data_0_995;
                  verilogPut_Key_2_973 <= verilogPut_Key_1_996;
                  verilogPut_Data_2_976 <= verilogPut_Data_1_999;
                  verilogPut_size_962 <= verilogPut_size_962 + 2;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                3: begin
                  verilogPut_Key_1_969 <= verilogPut_Key_0_992;
                  verilogPut_Data_1_972 <= verilogPut_Data_0_995;
                  verilogPut_Key_2_973 <= verilogPut_Key_1_996;
                  verilogPut_Data_2_976 <= verilogPut_Data_1_999;
                  verilogPut_Key_3_977 <= verilogPut_Key_2_1000;
                  verilogPut_Data_3_980 <= verilogPut_Data_2_1003;
                  verilogPut_size_962 <= verilogPut_size_962 + 3;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_989)
                0: begin
                  verilogPut_size_962 <= verilogPut_size_962 + 0;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                1: begin
                  verilogPut_Key_2_973 <= verilogPut_Key_0_992;
                  verilogPut_Data_2_976 <= verilogPut_Data_0_995;
                  verilogPut_size_962 <= verilogPut_size_962 + 1;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                2: begin
                  verilogPut_Key_2_973 <= verilogPut_Key_0_992;
                  verilogPut_Data_2_976 <= verilogPut_Data_0_995;
                  verilogPut_Key_3_977 <= verilogPut_Key_1_996;
                  verilogPut_Data_3_980 <= verilogPut_Data_1_999;
                  verilogPut_size_962 <= verilogPut_size_962 + 2;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_989)
                0: begin
                  verilogPut_size_962 <= verilogPut_size_962 + 0;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                1: begin
                  verilogPut_Key_3_977 <= verilogPut_Key_0_992;
                  verilogPut_Data_3_980 <= verilogPut_Data_0_995;
                  verilogPut_size_962 <= verilogPut_size_962 + 1;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_989)
                0: begin
                  verilogPut_size_962 <= verilogPut_size_962 + 0;
                  verilogPut_MergeSuccess_987 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        607: begin
          if (verilogPut_MergeSuccess_987 == 0) begin
            verilogPut_pc <= 627;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        608: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          verilogPut_success_1021 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        609: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_961;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_962;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_961;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_965;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_969;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_973;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_977;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_961;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_968;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_972;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_976;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_980;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        610: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        611: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        612: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        613: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        614: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        615: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        616: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        617: begin
          verilogPut_root_1024 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        618: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1024;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        619: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        620: begin
          verilogPut_next_1023 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1024;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1019;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1025 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        621: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1019;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1025;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        622: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        623: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1019;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1023;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        624: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        625: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        626: begin
          verilogPut_pc <= 627;
        end
        627: begin
          verilogPut_pc <= 628;
        end
        628: begin
          verilogPut_pc <= 629;
        end
        629: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 674;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        630: begin
          verilogPut_success_1086 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        631: begin
          verilogPut_size_1081 <= verilogPut_size_741;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        632: begin
          case (verilogPut_size_1081)
            1: begin
              verilogPut_indexLeft_1083 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1084 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_indexLeft_1083 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1084 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_indexLeft_1083 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1084 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        633: begin
          verilogPut_index_1026 <= verilogPut_indexLeft_1083;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        634: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1026;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1026;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1026;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1026;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        635: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        636: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        637: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        638: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        639: begin
          verilogPut_size_1027 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1028 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1030 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1033 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1034 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1037 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1038 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1041 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1042 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1045 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        640: begin
          verilogPut_index_1053 <= verilogPut_indexRight_1084;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        641: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1053;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1053;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1053;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1053;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        642: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        643: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        644: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        645: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        646: begin
          verilogPut_size_1054 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1055 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1057 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1060 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1061 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1064 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1065 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1068 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1069 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1072 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        647: begin
          if (verilogPut_isLeaf_1028 == 0) begin
            verilogPut_pc <= 649;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        648: begin
          verilogPut_pc <= 674;
        end
        649: begin
          if (verilogPut_isLeaf_1055 == 0) begin
            verilogPut_pc <= 651;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        650: begin
          verilogPut_pc <= 674;
        end
        651: begin
          case (verilogPut_size_741)
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            4: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_size_741 <= verilogPut_size_741-1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        652: begin
          verilogPut_MergeSuccess_1052 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        653: begin
          case (verilogPut_size_1027)
            0: begin
              case (verilogPut_size_1054)
                0: begin
                  verilogPut_Key_0_1030 <= verilogPut_Key_761;
                  verilogPut_Data_1_1037 <= verilogPut_Data_0_1060;
                  verilogPut_size_1027 <= verilogPut_size_1027 + 1;
                  verilogPut_MergeSuccess_1052 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1030 <= verilogPut_Key_761;
                  verilogPut_Key_1_1034 <= verilogPut_Key_0_1057;
                  verilogPut_Data_1_1037 <= verilogPut_Data_0_1060;
                  verilogPut_Data_2_1041 <= verilogPut_Data_1_1064;
                  verilogPut_size_1027 <= verilogPut_size_1027 + 2;
                  verilogPut_MergeSuccess_1052 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1030 <= verilogPut_Key_761;
                  verilogPut_Key_1_1034 <= verilogPut_Key_0_1057;
                  verilogPut_Data_1_1037 <= verilogPut_Data_0_1060;
                  verilogPut_Key_2_1038 <= verilogPut_Key_1_1061;
                  verilogPut_Data_2_1041 <= verilogPut_Data_1_1064;
                  verilogPut_Data_3_1045 <= verilogPut_Data_2_1068;
                  verilogPut_size_1027 <= verilogPut_size_1027 + 3;
                  verilogPut_MergeSuccess_1052 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1054)
                0: begin
                  verilogPut_Key_1_1034 <= verilogPut_Key_761;
                  verilogPut_Data_2_1041 <= verilogPut_Data_0_1060;
                  verilogPut_size_1027 <= verilogPut_size_1027 + 1;
                  verilogPut_MergeSuccess_1052 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1034 <= verilogPut_Key_761;
                  verilogPut_Key_2_1038 <= verilogPut_Key_0_1057;
                  verilogPut_Data_2_1041 <= verilogPut_Data_0_1060;
                  verilogPut_Data_3_1045 <= verilogPut_Data_1_1064;
                  verilogPut_size_1027 <= verilogPut_size_1027 + 2;
                  verilogPut_MergeSuccess_1052 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1054)
                0: begin
                  verilogPut_Key_2_1038 <= verilogPut_Key_761;
                  verilogPut_Data_3_1045 <= verilogPut_Data_0_1060;
                  verilogPut_size_1027 <= verilogPut_size_1027 + 1;
                  verilogPut_MergeSuccess_1052 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1054)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1054)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        654: begin
          if (verilogPut_MergeSuccess_1052 == 0) begin
            verilogPut_pc <= 674;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        655: begin
          verilogPut_success_1086 <= 1;
          case (verilogPut_size_741)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1083;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1083;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1083;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1083;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        656: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1026;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1027;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1026;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1030;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1034;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1038;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1042;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1026;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1033;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1037;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1041;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1045;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        657: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        658: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        659: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        660: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        661: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        662: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        663: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        664: begin
          verilogPut_root_1089 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        665: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1089;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        666: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        667: begin
          verilogPut_next_1088 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1089;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1084;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1090 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        668: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1084;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1090;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        669: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        670: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1084;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1088;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        671: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        672: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        673: begin
          verilogPut_pc <= 674;
        end
        674: begin
          verilogPut_index_740 <= verilogPut_position_767;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        675: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        676: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        677: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        678: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        679: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        680: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        681: begin
          verilogPut_index_768 <= 2;
          verilogPut_within_769 <= verilogPut_size_741>=3 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        682: begin
          if (verilogPut_within_769 == 0) begin
            verilogPut_pc <= 775;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        683: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 727;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        684: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_indexLeft_1147 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1148 <= verilogPut_Data_1_751;
            end
            1: begin
              verilogPut_indexLeft_1147 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1148 <= verilogPut_Data_2_755;
            end
            2: begin
              verilogPut_indexLeft_1147 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1148 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        685: begin
          verilogPut_index_1091 <= verilogPut_indexLeft_1147;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        686: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1091;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1091;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1091;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1091;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        687: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        688: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        689: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        690: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        691: begin
          verilogPut_size_1092 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1093 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1095 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1098 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1099 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1102 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1103 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1106 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1107 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1110 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        692: begin
          verilogPut_index_1118 <= verilogPut_indexRight_1148;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        693: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1118;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1118;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1118;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1118;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        694: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        695: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        696: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        697: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        698: begin
          verilogPut_size_1119 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1120 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1122 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1125 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1126 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1129 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1130 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1133 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1134 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1137 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        699: begin
          if (verilogPut_isLeaf_1093 == 0) begin
            verilogPut_pc <= 727;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        700: begin
          if (verilogPut_isLeaf_1120 == 0) begin
            verilogPut_pc <= 726;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        701: begin
          verilogPut_MergeSuccess_1117 <= 0;
          case (verilogPut_size_1092)
            0: begin
              case (verilogPut_size_1119)
                0: begin
                  verilogPut_size_1092 <= verilogPut_size_1092 + 0;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1095 <= verilogPut_Key_0_1122;
                  verilogPut_Data_0_1098 <= verilogPut_Data_0_1125;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 1;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1095 <= verilogPut_Key_0_1122;
                  verilogPut_Data_0_1098 <= verilogPut_Data_0_1125;
                  verilogPut_Key_1_1099 <= verilogPut_Key_1_1126;
                  verilogPut_Data_1_1102 <= verilogPut_Data_1_1129;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 2;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                3: begin
                  verilogPut_Key_0_1095 <= verilogPut_Key_0_1122;
                  verilogPut_Data_0_1098 <= verilogPut_Data_0_1125;
                  verilogPut_Key_1_1099 <= verilogPut_Key_1_1126;
                  verilogPut_Data_1_1102 <= verilogPut_Data_1_1129;
                  verilogPut_Key_2_1103 <= verilogPut_Key_2_1130;
                  verilogPut_Data_2_1106 <= verilogPut_Data_2_1133;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 3;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                4: begin
                  verilogPut_Key_0_1095 <= verilogPut_Key_0_1122;
                  verilogPut_Data_0_1098 <= verilogPut_Data_0_1125;
                  verilogPut_Key_1_1099 <= verilogPut_Key_1_1126;
                  verilogPut_Data_1_1102 <= verilogPut_Data_1_1129;
                  verilogPut_Key_2_1103 <= verilogPut_Key_2_1130;
                  verilogPut_Data_2_1106 <= verilogPut_Data_2_1133;
                  verilogPut_Key_3_1107 <= verilogPut_Key_3_1134;
                  verilogPut_Data_3_1110 <= verilogPut_Data_3_1137;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 4;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1119)
                0: begin
                  verilogPut_size_1092 <= verilogPut_size_1092 + 0;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1099 <= verilogPut_Key_0_1122;
                  verilogPut_Data_1_1102 <= verilogPut_Data_0_1125;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 1;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                2: begin
                  verilogPut_Key_1_1099 <= verilogPut_Key_0_1122;
                  verilogPut_Data_1_1102 <= verilogPut_Data_0_1125;
                  verilogPut_Key_2_1103 <= verilogPut_Key_1_1126;
                  verilogPut_Data_2_1106 <= verilogPut_Data_1_1129;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 2;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                3: begin
                  verilogPut_Key_1_1099 <= verilogPut_Key_0_1122;
                  verilogPut_Data_1_1102 <= verilogPut_Data_0_1125;
                  verilogPut_Key_2_1103 <= verilogPut_Key_1_1126;
                  verilogPut_Data_2_1106 <= verilogPut_Data_1_1129;
                  verilogPut_Key_3_1107 <= verilogPut_Key_2_1130;
                  verilogPut_Data_3_1110 <= verilogPut_Data_2_1133;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 3;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1119)
                0: begin
                  verilogPut_size_1092 <= verilogPut_size_1092 + 0;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                1: begin
                  verilogPut_Key_2_1103 <= verilogPut_Key_0_1122;
                  verilogPut_Data_2_1106 <= verilogPut_Data_0_1125;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 1;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                2: begin
                  verilogPut_Key_2_1103 <= verilogPut_Key_0_1122;
                  verilogPut_Data_2_1106 <= verilogPut_Data_0_1125;
                  verilogPut_Key_3_1107 <= verilogPut_Key_1_1126;
                  verilogPut_Data_3_1110 <= verilogPut_Data_1_1129;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 2;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1119)
                0: begin
                  verilogPut_size_1092 <= verilogPut_size_1092 + 0;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                1: begin
                  verilogPut_Key_3_1107 <= verilogPut_Key_0_1122;
                  verilogPut_Data_3_1110 <= verilogPut_Data_0_1125;
                  verilogPut_size_1092 <= verilogPut_size_1092 + 1;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1119)
                0: begin
                  verilogPut_size_1092 <= verilogPut_size_1092 + 0;
                  verilogPut_MergeSuccess_1117 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        702: begin
          if (verilogPut_MergeSuccess_1117 == 0) begin
            verilogPut_pc <= 725;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        703: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          if (0>= verilogPut_index_768) begin
            verilogPut_Key_0_744 <= verilogPut_Key_1_748;
            verilogPut_Data_0_747 <= verilogPut_Data_1_751;
          end
          if (1>= verilogPut_index_768) begin
            verilogPut_Key_1_748 <= verilogPut_Key_2_752;
            verilogPut_Data_1_751 <= verilogPut_Data_2_755;
          end
          if (2>= verilogPut_index_768) begin
            verilogPut_Key_2_752 <= verilogPut_Key_3_756;
            verilogPut_Data_2_755 <= verilogPut_Data_3_759;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        704: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        705: begin
          if (verilogPut_index_768 == verilogPut_size_741) begin
            verilogPut_size_741 <= verilogPut_size_741+1;
          end
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1147;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1147;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1147;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1147;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        706: begin
          verilogPut_success_1150 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        707: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1091;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1092;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1091;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1095;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1099;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1103;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1107;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1091;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1098;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1102;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1106;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1110;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        708: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        709: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        710: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        711: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        712: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        713: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        714: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        715: begin
          verilogPut_root_1153 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        716: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1153;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        717: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        718: begin
          verilogPut_next_1152 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1153;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1148;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1154 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        719: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1148;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1154;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        720: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        721: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1148;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1152;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        722: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        723: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        724: begin
          verilogPut_pc <= 725;
        end
        725: begin
          verilogPut_pc <= 726;
        end
        726: begin
          verilogPut_pc <= 727;
        end
        727: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 774;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        728: begin
          verilogPut_success_1216 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        729: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_indexLeft_1213 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1214 <= verilogPut_Data_1_751;
            end
            1: begin
              verilogPut_indexLeft_1213 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1214 <= verilogPut_Data_2_755;
            end
            2: begin
              verilogPut_indexLeft_1213 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1214 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        730: begin
          verilogPut_index_1155 <= verilogPut_indexLeft_1213;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        731: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1155;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1155;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1155;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1155;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        732: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        733: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        734: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        735: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        736: begin
          verilogPut_size_1156 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1157 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1159 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1162 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1163 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1166 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1167 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1170 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1171 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1174 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        737: begin
          verilogPut_index_1182 <= verilogPut_indexRight_1214;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        738: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1182;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1182;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1182;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1182;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        739: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        740: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        741: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        742: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        743: begin
          verilogPut_size_1183 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1184 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1186 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1189 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1190 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1193 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1194 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1197 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1198 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1201 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        744: begin
          if (verilogPut_isLeaf_1157 == 0) begin
            verilogPut_pc <= 746;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        745: begin
          verilogPut_pc <= 774;
        end
        746: begin
          if (verilogPut_isLeaf_1184 == 0) begin
            verilogPut_pc <= 748;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        747: begin
          verilogPut_pc <= 774;
        end
        748: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_midKey_1215 <= verilogPut_Key_0_744;
            end
            1: begin
              verilogPut_midKey_1215 <= verilogPut_Key_1_748;
            end
            2: begin
              verilogPut_midKey_1215 <= verilogPut_Key_2_752;
            end
            3: begin
              verilogPut_midKey_1215 <= verilogPut_Key_3_756;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        749: begin
          verilogPut_MergeSuccess_1181 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        750: begin
          case (verilogPut_size_1156)
            0: begin
              case (verilogPut_size_1183)
                0: begin
                  verilogPut_Key_0_1159 <= verilogPut_midKey_1215;
                  verilogPut_Data_1_1166 <= verilogPut_Data_0_1189;
                  verilogPut_size_1156 <= verilogPut_size_1156 + 1;
                  verilogPut_MergeSuccess_1181 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1159 <= verilogPut_midKey_1215;
                  verilogPut_Key_1_1163 <= verilogPut_Key_0_1186;
                  verilogPut_Data_1_1166 <= verilogPut_Data_0_1189;
                  verilogPut_Data_2_1170 <= verilogPut_Data_1_1193;
                  verilogPut_size_1156 <= verilogPut_size_1156 + 2;
                  verilogPut_MergeSuccess_1181 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1159 <= verilogPut_midKey_1215;
                  verilogPut_Key_1_1163 <= verilogPut_Key_0_1186;
                  verilogPut_Data_1_1166 <= verilogPut_Data_0_1189;
                  verilogPut_Key_2_1167 <= verilogPut_Key_1_1190;
                  verilogPut_Data_2_1170 <= verilogPut_Data_1_1193;
                  verilogPut_Data_3_1174 <= verilogPut_Data_2_1197;
                  verilogPut_size_1156 <= verilogPut_size_1156 + 3;
                  verilogPut_MergeSuccess_1181 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1183)
                0: begin
                  verilogPut_Key_1_1163 <= verilogPut_midKey_1215;
                  verilogPut_Data_2_1170 <= verilogPut_Data_0_1189;
                  verilogPut_size_1156 <= verilogPut_size_1156 + 1;
                  verilogPut_MergeSuccess_1181 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1163 <= verilogPut_midKey_1215;
                  verilogPut_Key_2_1167 <= verilogPut_Key_0_1186;
                  verilogPut_Data_2_1170 <= verilogPut_Data_0_1189;
                  verilogPut_Data_3_1174 <= verilogPut_Data_1_1193;
                  verilogPut_size_1156 <= verilogPut_size_1156 + 2;
                  verilogPut_MergeSuccess_1181 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1183)
                0: begin
                  verilogPut_Key_2_1167 <= verilogPut_midKey_1215;
                  verilogPut_Data_3_1174 <= verilogPut_Data_0_1189;
                  verilogPut_size_1156 <= verilogPut_size_1156 + 1;
                  verilogPut_MergeSuccess_1181 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1183)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1183)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        751: begin
          if (verilogPut_MergeSuccess_1181 == 0) begin
            verilogPut_pc <= 774;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        752: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          if (0>= verilogPut_index_768) begin
            verilogPut_Key_0_744 <= verilogPut_Key_1_748;
            verilogPut_Data_0_747 <= verilogPut_Data_1_751;
          end
          if (1>= verilogPut_index_768) begin
            verilogPut_Key_1_748 <= verilogPut_Key_2_752;
            verilogPut_Data_1_751 <= verilogPut_Data_2_755;
          end
          if (2>= verilogPut_index_768) begin
            verilogPut_Key_2_752 <= verilogPut_Key_3_756;
            verilogPut_Data_2_755 <= verilogPut_Data_3_759;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        753: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        754: begin
          if (verilogPut_index_768 == verilogPut_size_741) begin
            verilogPut_size_741 <= verilogPut_size_741+1;
          end
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1213;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1213;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1213;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1213;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        755: begin
          verilogPut_success_1216 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        756: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1155;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1156;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1155;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1159;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1163;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1167;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1171;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1155;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1162;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1166;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1170;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1174;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        757: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        758: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        759: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        760: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        761: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        762: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        763: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        764: begin
          verilogPut_root_1219 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        765: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1219;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        766: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        767: begin
          verilogPut_next_1218 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1219;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1214;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1220 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        768: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1214;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1220;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        769: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        770: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1214;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1218;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        771: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        772: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        773: begin
          verilogPut_pc <= 774;
        end
        774: begin
          verilogPut_pc <= 775;
        end
        775: begin
          verilogPut_index_740 <= verilogPut_position_767;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        776: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        777: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        778: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        779: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        780: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        781: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        782: begin
          verilogPut_index_768 <= 1;
          verilogPut_within_769 <= verilogPut_size_741>=2 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        783: begin
          if (verilogPut_within_769 == 0) begin
            verilogPut_pc <= 876;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        784: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 828;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        785: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_indexLeft_1277 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1278 <= verilogPut_Data_1_751;
            end
            1: begin
              verilogPut_indexLeft_1277 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1278 <= verilogPut_Data_2_755;
            end
            2: begin
              verilogPut_indexLeft_1277 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1278 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        786: begin
          verilogPut_index_1221 <= verilogPut_indexLeft_1277;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        787: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1221;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1221;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1221;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1221;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        788: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        789: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        790: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        791: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        792: begin
          verilogPut_size_1222 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1223 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1225 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1228 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1229 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1232 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1233 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1236 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1237 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1240 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        793: begin
          verilogPut_index_1248 <= verilogPut_indexRight_1278;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        794: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1248;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1248;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1248;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1248;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        795: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        796: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        797: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        798: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        799: begin
          verilogPut_size_1249 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1250 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1252 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1255 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1256 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1259 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1260 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1263 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1264 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1267 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        800: begin
          if (verilogPut_isLeaf_1223 == 0) begin
            verilogPut_pc <= 828;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        801: begin
          if (verilogPut_isLeaf_1250 == 0) begin
            verilogPut_pc <= 827;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        802: begin
          verilogPut_MergeSuccess_1247 <= 0;
          case (verilogPut_size_1222)
            0: begin
              case (verilogPut_size_1249)
                0: begin
                  verilogPut_size_1222 <= verilogPut_size_1222 + 0;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1225 <= verilogPut_Key_0_1252;
                  verilogPut_Data_0_1228 <= verilogPut_Data_0_1255;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 1;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1225 <= verilogPut_Key_0_1252;
                  verilogPut_Data_0_1228 <= verilogPut_Data_0_1255;
                  verilogPut_Key_1_1229 <= verilogPut_Key_1_1256;
                  verilogPut_Data_1_1232 <= verilogPut_Data_1_1259;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 2;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                3: begin
                  verilogPut_Key_0_1225 <= verilogPut_Key_0_1252;
                  verilogPut_Data_0_1228 <= verilogPut_Data_0_1255;
                  verilogPut_Key_1_1229 <= verilogPut_Key_1_1256;
                  verilogPut_Data_1_1232 <= verilogPut_Data_1_1259;
                  verilogPut_Key_2_1233 <= verilogPut_Key_2_1260;
                  verilogPut_Data_2_1236 <= verilogPut_Data_2_1263;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 3;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                4: begin
                  verilogPut_Key_0_1225 <= verilogPut_Key_0_1252;
                  verilogPut_Data_0_1228 <= verilogPut_Data_0_1255;
                  verilogPut_Key_1_1229 <= verilogPut_Key_1_1256;
                  verilogPut_Data_1_1232 <= verilogPut_Data_1_1259;
                  verilogPut_Key_2_1233 <= verilogPut_Key_2_1260;
                  verilogPut_Data_2_1236 <= verilogPut_Data_2_1263;
                  verilogPut_Key_3_1237 <= verilogPut_Key_3_1264;
                  verilogPut_Data_3_1240 <= verilogPut_Data_3_1267;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 4;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1249)
                0: begin
                  verilogPut_size_1222 <= verilogPut_size_1222 + 0;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1229 <= verilogPut_Key_0_1252;
                  verilogPut_Data_1_1232 <= verilogPut_Data_0_1255;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 1;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                2: begin
                  verilogPut_Key_1_1229 <= verilogPut_Key_0_1252;
                  verilogPut_Data_1_1232 <= verilogPut_Data_0_1255;
                  verilogPut_Key_2_1233 <= verilogPut_Key_1_1256;
                  verilogPut_Data_2_1236 <= verilogPut_Data_1_1259;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 2;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                3: begin
                  verilogPut_Key_1_1229 <= verilogPut_Key_0_1252;
                  verilogPut_Data_1_1232 <= verilogPut_Data_0_1255;
                  verilogPut_Key_2_1233 <= verilogPut_Key_1_1256;
                  verilogPut_Data_2_1236 <= verilogPut_Data_1_1259;
                  verilogPut_Key_3_1237 <= verilogPut_Key_2_1260;
                  verilogPut_Data_3_1240 <= verilogPut_Data_2_1263;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 3;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1249)
                0: begin
                  verilogPut_size_1222 <= verilogPut_size_1222 + 0;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                1: begin
                  verilogPut_Key_2_1233 <= verilogPut_Key_0_1252;
                  verilogPut_Data_2_1236 <= verilogPut_Data_0_1255;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 1;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                2: begin
                  verilogPut_Key_2_1233 <= verilogPut_Key_0_1252;
                  verilogPut_Data_2_1236 <= verilogPut_Data_0_1255;
                  verilogPut_Key_3_1237 <= verilogPut_Key_1_1256;
                  verilogPut_Data_3_1240 <= verilogPut_Data_1_1259;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 2;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1249)
                0: begin
                  verilogPut_size_1222 <= verilogPut_size_1222 + 0;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                1: begin
                  verilogPut_Key_3_1237 <= verilogPut_Key_0_1252;
                  verilogPut_Data_3_1240 <= verilogPut_Data_0_1255;
                  verilogPut_size_1222 <= verilogPut_size_1222 + 1;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1249)
                0: begin
                  verilogPut_size_1222 <= verilogPut_size_1222 + 0;
                  verilogPut_MergeSuccess_1247 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        803: begin
          if (verilogPut_MergeSuccess_1247 == 0) begin
            verilogPut_pc <= 826;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        804: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          if (0>= verilogPut_index_768) begin
            verilogPut_Key_0_744 <= verilogPut_Key_1_748;
            verilogPut_Data_0_747 <= verilogPut_Data_1_751;
          end
          if (1>= verilogPut_index_768) begin
            verilogPut_Key_1_748 <= verilogPut_Key_2_752;
            verilogPut_Data_1_751 <= verilogPut_Data_2_755;
          end
          if (2>= verilogPut_index_768) begin
            verilogPut_Key_2_752 <= verilogPut_Key_3_756;
            verilogPut_Data_2_755 <= verilogPut_Data_3_759;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        805: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        806: begin
          if (verilogPut_index_768 == verilogPut_size_741) begin
            verilogPut_size_741 <= verilogPut_size_741+1;
          end
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1277;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1277;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1277;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1277;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        807: begin
          verilogPut_success_1280 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        808: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1221;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1222;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1221;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1225;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1229;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1233;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1237;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1221;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1228;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1232;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1236;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1240;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        809: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        810: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        811: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        812: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        813: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        814: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        815: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        816: begin
          verilogPut_root_1283 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        817: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1283;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        818: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        819: begin
          verilogPut_next_1282 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1283;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1278;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1284 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        820: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1278;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1284;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        821: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        822: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1278;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1282;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        823: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        824: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        825: begin
          verilogPut_pc <= 826;
        end
        826: begin
          verilogPut_pc <= 827;
        end
        827: begin
          verilogPut_pc <= 828;
        end
        828: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 875;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        829: begin
          verilogPut_success_1346 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        830: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_indexLeft_1343 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1344 <= verilogPut_Data_1_751;
            end
            1: begin
              verilogPut_indexLeft_1343 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1344 <= verilogPut_Data_2_755;
            end
            2: begin
              verilogPut_indexLeft_1343 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1344 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        831: begin
          verilogPut_index_1285 <= verilogPut_indexLeft_1343;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        832: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1285;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1285;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1285;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1285;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        833: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        834: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        835: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        836: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        837: begin
          verilogPut_size_1286 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1287 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1289 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1292 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1293 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1296 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1297 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1300 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1301 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1304 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        838: begin
          verilogPut_index_1312 <= verilogPut_indexRight_1344;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        839: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1312;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1312;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1312;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1312;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        840: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        841: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        842: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        843: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        844: begin
          verilogPut_size_1313 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1314 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1316 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1319 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1320 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1323 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1324 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1327 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1328 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1331 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        845: begin
          if (verilogPut_isLeaf_1287 == 0) begin
            verilogPut_pc <= 847;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        846: begin
          verilogPut_pc <= 875;
        end
        847: begin
          if (verilogPut_isLeaf_1314 == 0) begin
            verilogPut_pc <= 849;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        848: begin
          verilogPut_pc <= 875;
        end
        849: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_midKey_1345 <= verilogPut_Key_0_744;
            end
            1: begin
              verilogPut_midKey_1345 <= verilogPut_Key_1_748;
            end
            2: begin
              verilogPut_midKey_1345 <= verilogPut_Key_2_752;
            end
            3: begin
              verilogPut_midKey_1345 <= verilogPut_Key_3_756;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        850: begin
          verilogPut_MergeSuccess_1311 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        851: begin
          case (verilogPut_size_1286)
            0: begin
              case (verilogPut_size_1313)
                0: begin
                  verilogPut_Key_0_1289 <= verilogPut_midKey_1345;
                  verilogPut_Data_1_1296 <= verilogPut_Data_0_1319;
                  verilogPut_size_1286 <= verilogPut_size_1286 + 1;
                  verilogPut_MergeSuccess_1311 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1289 <= verilogPut_midKey_1345;
                  verilogPut_Key_1_1293 <= verilogPut_Key_0_1316;
                  verilogPut_Data_1_1296 <= verilogPut_Data_0_1319;
                  verilogPut_Data_2_1300 <= verilogPut_Data_1_1323;
                  verilogPut_size_1286 <= verilogPut_size_1286 + 2;
                  verilogPut_MergeSuccess_1311 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1289 <= verilogPut_midKey_1345;
                  verilogPut_Key_1_1293 <= verilogPut_Key_0_1316;
                  verilogPut_Data_1_1296 <= verilogPut_Data_0_1319;
                  verilogPut_Key_2_1297 <= verilogPut_Key_1_1320;
                  verilogPut_Data_2_1300 <= verilogPut_Data_1_1323;
                  verilogPut_Data_3_1304 <= verilogPut_Data_2_1327;
                  verilogPut_size_1286 <= verilogPut_size_1286 + 3;
                  verilogPut_MergeSuccess_1311 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1313)
                0: begin
                  verilogPut_Key_1_1293 <= verilogPut_midKey_1345;
                  verilogPut_Data_2_1300 <= verilogPut_Data_0_1319;
                  verilogPut_size_1286 <= verilogPut_size_1286 + 1;
                  verilogPut_MergeSuccess_1311 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1293 <= verilogPut_midKey_1345;
                  verilogPut_Key_2_1297 <= verilogPut_Key_0_1316;
                  verilogPut_Data_2_1300 <= verilogPut_Data_0_1319;
                  verilogPut_Data_3_1304 <= verilogPut_Data_1_1323;
                  verilogPut_size_1286 <= verilogPut_size_1286 + 2;
                  verilogPut_MergeSuccess_1311 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1313)
                0: begin
                  verilogPut_Key_2_1297 <= verilogPut_midKey_1345;
                  verilogPut_Data_3_1304 <= verilogPut_Data_0_1319;
                  verilogPut_size_1286 <= verilogPut_size_1286 + 1;
                  verilogPut_MergeSuccess_1311 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1313)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1313)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        852: begin
          if (verilogPut_MergeSuccess_1311 == 0) begin
            verilogPut_pc <= 875;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        853: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          if (0>= verilogPut_index_768) begin
            verilogPut_Key_0_744 <= verilogPut_Key_1_748;
            verilogPut_Data_0_747 <= verilogPut_Data_1_751;
          end
          if (1>= verilogPut_index_768) begin
            verilogPut_Key_1_748 <= verilogPut_Key_2_752;
            verilogPut_Data_1_751 <= verilogPut_Data_2_755;
          end
          if (2>= verilogPut_index_768) begin
            verilogPut_Key_2_752 <= verilogPut_Key_3_756;
            verilogPut_Data_2_755 <= verilogPut_Data_3_759;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        854: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        855: begin
          if (verilogPut_index_768 == verilogPut_size_741) begin
            verilogPut_size_741 <= verilogPut_size_741+1;
          end
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1343;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1343;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1343;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1343;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        856: begin
          verilogPut_success_1346 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        857: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1285;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1286;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1285;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1289;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1293;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1297;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1301;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1285;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1292;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1296;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1300;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1304;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        858: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        859: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        860: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        861: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        862: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        863: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        864: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        865: begin
          verilogPut_root_1349 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        866: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1349;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        867: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        868: begin
          verilogPut_next_1348 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1349;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1344;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1350 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        869: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1344;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1350;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        870: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        871: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1344;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1348;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        872: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        873: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        874: begin
          verilogPut_pc <= 875;
        end
        875: begin
          verilogPut_pc <= 876;
        end
        876: begin
          verilogPut_index_740 <= verilogPut_position_767;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        877: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        878: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        879: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        880: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        881: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        882: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        883: begin
          verilogPut_index_768 <= 0;
          verilogPut_within_769 <= verilogPut_size_741>=1 ? 1 : 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        884: begin
          if (verilogPut_within_769 == 0) begin
            verilogPut_pc <= 977;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        885: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 929;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        886: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_indexLeft_1407 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1408 <= verilogPut_Data_1_751;
            end
            1: begin
              verilogPut_indexLeft_1407 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1408 <= verilogPut_Data_2_755;
            end
            2: begin
              verilogPut_indexLeft_1407 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1408 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        887: begin
          verilogPut_index_1351 <= verilogPut_indexLeft_1407;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        888: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1351;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1351;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1351;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1351;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        889: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        890: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        891: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        892: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        893: begin
          verilogPut_size_1352 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1353 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1355 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1358 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1359 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1362 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1363 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1366 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1367 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1370 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        894: begin
          verilogPut_index_1378 <= verilogPut_indexRight_1408;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        895: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1378;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1378;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1378;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1378;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        896: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        897: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        898: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        899: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        900: begin
          verilogPut_size_1379 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1380 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1382 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1385 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1386 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1389 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1390 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1393 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1394 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1397 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        901: begin
          if (verilogPut_isLeaf_1353 == 0) begin
            verilogPut_pc <= 929;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        902: begin
          if (verilogPut_isLeaf_1380 == 0) begin
            verilogPut_pc <= 928;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        903: begin
          verilogPut_MergeSuccess_1377 <= 0;
          case (verilogPut_size_1352)
            0: begin
              case (verilogPut_size_1379)
                0: begin
                  verilogPut_size_1352 <= verilogPut_size_1352 + 0;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1355 <= verilogPut_Key_0_1382;
                  verilogPut_Data_0_1358 <= verilogPut_Data_0_1385;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 1;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1355 <= verilogPut_Key_0_1382;
                  verilogPut_Data_0_1358 <= verilogPut_Data_0_1385;
                  verilogPut_Key_1_1359 <= verilogPut_Key_1_1386;
                  verilogPut_Data_1_1362 <= verilogPut_Data_1_1389;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 2;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                3: begin
                  verilogPut_Key_0_1355 <= verilogPut_Key_0_1382;
                  verilogPut_Data_0_1358 <= verilogPut_Data_0_1385;
                  verilogPut_Key_1_1359 <= verilogPut_Key_1_1386;
                  verilogPut_Data_1_1362 <= verilogPut_Data_1_1389;
                  verilogPut_Key_2_1363 <= verilogPut_Key_2_1390;
                  verilogPut_Data_2_1366 <= verilogPut_Data_2_1393;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 3;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                4: begin
                  verilogPut_Key_0_1355 <= verilogPut_Key_0_1382;
                  verilogPut_Data_0_1358 <= verilogPut_Data_0_1385;
                  verilogPut_Key_1_1359 <= verilogPut_Key_1_1386;
                  verilogPut_Data_1_1362 <= verilogPut_Data_1_1389;
                  verilogPut_Key_2_1363 <= verilogPut_Key_2_1390;
                  verilogPut_Data_2_1366 <= verilogPut_Data_2_1393;
                  verilogPut_Key_3_1367 <= verilogPut_Key_3_1394;
                  verilogPut_Data_3_1370 <= verilogPut_Data_3_1397;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 4;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1379)
                0: begin
                  verilogPut_size_1352 <= verilogPut_size_1352 + 0;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1359 <= verilogPut_Key_0_1382;
                  verilogPut_Data_1_1362 <= verilogPut_Data_0_1385;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 1;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                2: begin
                  verilogPut_Key_1_1359 <= verilogPut_Key_0_1382;
                  verilogPut_Data_1_1362 <= verilogPut_Data_0_1385;
                  verilogPut_Key_2_1363 <= verilogPut_Key_1_1386;
                  verilogPut_Data_2_1366 <= verilogPut_Data_1_1389;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 2;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                3: begin
                  verilogPut_Key_1_1359 <= verilogPut_Key_0_1382;
                  verilogPut_Data_1_1362 <= verilogPut_Data_0_1385;
                  verilogPut_Key_2_1363 <= verilogPut_Key_1_1386;
                  verilogPut_Data_2_1366 <= verilogPut_Data_1_1389;
                  verilogPut_Key_3_1367 <= verilogPut_Key_2_1390;
                  verilogPut_Data_3_1370 <= verilogPut_Data_2_1393;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 3;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1379)
                0: begin
                  verilogPut_size_1352 <= verilogPut_size_1352 + 0;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                1: begin
                  verilogPut_Key_2_1363 <= verilogPut_Key_0_1382;
                  verilogPut_Data_2_1366 <= verilogPut_Data_0_1385;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 1;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                2: begin
                  verilogPut_Key_2_1363 <= verilogPut_Key_0_1382;
                  verilogPut_Data_2_1366 <= verilogPut_Data_0_1385;
                  verilogPut_Key_3_1367 <= verilogPut_Key_1_1386;
                  verilogPut_Data_3_1370 <= verilogPut_Data_1_1389;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 2;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1379)
                0: begin
                  verilogPut_size_1352 <= verilogPut_size_1352 + 0;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                1: begin
                  verilogPut_Key_3_1367 <= verilogPut_Key_0_1382;
                  verilogPut_Data_3_1370 <= verilogPut_Data_0_1385;
                  verilogPut_size_1352 <= verilogPut_size_1352 + 1;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1379)
                0: begin
                  verilogPut_size_1352 <= verilogPut_size_1352 + 0;
                  verilogPut_MergeSuccess_1377 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        904: begin
          if (verilogPut_MergeSuccess_1377 == 0) begin
            verilogPut_pc <= 927;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        905: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          if (0>= verilogPut_index_768) begin
            verilogPut_Key_0_744 <= verilogPut_Key_1_748;
            verilogPut_Data_0_747 <= verilogPut_Data_1_751;
          end
          if (1>= verilogPut_index_768) begin
            verilogPut_Key_1_748 <= verilogPut_Key_2_752;
            verilogPut_Data_1_751 <= verilogPut_Data_2_755;
          end
          if (2>= verilogPut_index_768) begin
            verilogPut_Key_2_752 <= verilogPut_Key_3_756;
            verilogPut_Data_2_755 <= verilogPut_Data_3_759;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        906: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        907: begin
          if (verilogPut_index_768 == verilogPut_size_741) begin
            verilogPut_size_741 <= verilogPut_size_741+1;
          end
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1407;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1407;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1407;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1407;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        908: begin
          verilogPut_success_1410 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        909: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1351;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1352;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1351;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1355;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1359;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1363;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1367;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1351;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1358;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1362;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1366;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1370;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        910: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        911: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        912: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        913: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        914: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        915: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        916: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        917: begin
          verilogPut_root_1413 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        918: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1413;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        919: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        920: begin
          verilogPut_next_1412 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1413;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1408;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1414 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        921: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1408;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1414;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        922: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        923: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1408;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1412;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        924: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        925: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        926: begin
          verilogPut_pc <= 927;
        end
        927: begin
          verilogPut_pc <= 928;
        end
        928: begin
          verilogPut_pc <= 929;
        end
        929: begin
          if (verilogPut_position_767 == 0 && verilogPut_size_741 > 1) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
          else begin
            if (verilogPut_position_767 == 0 || verilogPut_size_741 < 1) begin
              verilogPut_pc <= 976;
            end
            else begin
              verilogPut_pc <= verilogPut_pc + 1;
            end
          end
        end
        930: begin
          verilogPut_success_1476 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        931: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_indexLeft_1473 <= verilogPut_Data_0_747;
              verilogPut_indexRight_1474 <= verilogPut_Data_1_751;
            end
            1: begin
              verilogPut_indexLeft_1473 <= verilogPut_Data_1_751;
              verilogPut_indexRight_1474 <= verilogPut_Data_2_755;
            end
            2: begin
              verilogPut_indexLeft_1473 <= verilogPut_Data_2_755;
              verilogPut_indexRight_1474 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        932: begin
          verilogPut_index_1415 <= verilogPut_indexLeft_1473;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        933: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1415;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1415;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1415;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1415;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        934: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        935: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        936: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        937: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        938: begin
          verilogPut_size_1416 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1417 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1419 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1422 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1423 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1426 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1427 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1430 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1431 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1434 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        939: begin
          verilogPut_index_1442 <= verilogPut_indexRight_1474;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        940: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_1442;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_1442;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_1442;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_1442;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        941: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        942: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        943: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        944: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        945: begin
          verilogPut_size_1443 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_1444 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_1446 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_1449 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_1450 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_1453 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_1454 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_1457 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_1458 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_1461 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        946: begin
          if (verilogPut_isLeaf_1417 == 0) begin
            verilogPut_pc <= 948;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        947: begin
          verilogPut_pc <= 976;
        end
        948: begin
          if (verilogPut_isLeaf_1444 == 0) begin
            verilogPut_pc <= 950;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        949: begin
          verilogPut_pc <= 976;
        end
        950: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_midKey_1475 <= verilogPut_Key_0_744;
            end
            1: begin
              verilogPut_midKey_1475 <= verilogPut_Key_1_748;
            end
            2: begin
              verilogPut_midKey_1475 <= verilogPut_Key_2_752;
            end
            3: begin
              verilogPut_midKey_1475 <= verilogPut_Key_3_756;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        951: begin
          verilogPut_MergeSuccess_1441 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        952: begin
          case (verilogPut_size_1416)
            0: begin
              case (verilogPut_size_1443)
                0: begin
                  verilogPut_Key_0_1419 <= verilogPut_midKey_1475;
                  verilogPut_Data_1_1426 <= verilogPut_Data_0_1449;
                  verilogPut_size_1416 <= verilogPut_size_1416 + 1;
                  verilogPut_MergeSuccess_1441 <= 1;
                end
                1: begin
                  verilogPut_Key_0_1419 <= verilogPut_midKey_1475;
                  verilogPut_Key_1_1423 <= verilogPut_Key_0_1446;
                  verilogPut_Data_1_1426 <= verilogPut_Data_0_1449;
                  verilogPut_Data_2_1430 <= verilogPut_Data_1_1453;
                  verilogPut_size_1416 <= verilogPut_size_1416 + 2;
                  verilogPut_MergeSuccess_1441 <= 1;
                end
                2: begin
                  verilogPut_Key_0_1419 <= verilogPut_midKey_1475;
                  verilogPut_Key_1_1423 <= verilogPut_Key_0_1446;
                  verilogPut_Data_1_1426 <= verilogPut_Data_0_1449;
                  verilogPut_Key_2_1427 <= verilogPut_Key_1_1450;
                  verilogPut_Data_2_1430 <= verilogPut_Data_1_1453;
                  verilogPut_Data_3_1434 <= verilogPut_Data_2_1457;
                  verilogPut_size_1416 <= verilogPut_size_1416 + 3;
                  verilogPut_MergeSuccess_1441 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (verilogPut_size_1443)
                0: begin
                  verilogPut_Key_1_1423 <= verilogPut_midKey_1475;
                  verilogPut_Data_2_1430 <= verilogPut_Data_0_1449;
                  verilogPut_size_1416 <= verilogPut_size_1416 + 1;
                  verilogPut_MergeSuccess_1441 <= 1;
                end
                1: begin
                  verilogPut_Key_1_1423 <= verilogPut_midKey_1475;
                  verilogPut_Key_2_1427 <= verilogPut_Key_0_1446;
                  verilogPut_Data_2_1430 <= verilogPut_Data_0_1449;
                  verilogPut_Data_3_1434 <= verilogPut_Data_1_1453;
                  verilogPut_size_1416 <= verilogPut_size_1416 + 2;
                  verilogPut_MergeSuccess_1441 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (verilogPut_size_1443)
                0: begin
                  verilogPut_Key_2_1427 <= verilogPut_midKey_1475;
                  verilogPut_Data_3_1434 <= verilogPut_Data_0_1449;
                  verilogPut_size_1416 <= verilogPut_size_1416 + 1;
                  verilogPut_MergeSuccess_1441 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (verilogPut_size_1443)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (verilogPut_size_1443)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        953: begin
          if (verilogPut_MergeSuccess_1441 == 0) begin
            verilogPut_pc <= 976;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        954: begin
          verilogPut_size_741 <= verilogPut_size_741-1;
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          if (0>= verilogPut_index_768) begin
            verilogPut_Key_0_744 <= verilogPut_Key_1_748;
            verilogPut_Data_0_747 <= verilogPut_Data_1_751;
          end
          if (1>= verilogPut_index_768) begin
            verilogPut_Key_1_748 <= verilogPut_Key_2_752;
            verilogPut_Data_1_751 <= verilogPut_Data_2_755;
          end
          if (2>= verilogPut_index_768) begin
            verilogPut_Key_2_752 <= verilogPut_Key_3_756;
            verilogPut_Data_2_755 <= verilogPut_Data_3_759;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        955: begin
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_761 <= verilogPut_Key_0_744;
              verilogPut_Data_763 <= verilogPut_Data_0_747;
            end
            1: begin
              verilogPut_Key_761 <= verilogPut_Key_1_748;
              verilogPut_Data_763 <= verilogPut_Data_1_751;
            end
            2: begin
              verilogPut_Key_761 <= verilogPut_Key_2_752;
              verilogPut_Data_763 <= verilogPut_Data_2_755;
            end
            3: begin
              verilogPut_Key_761 <= verilogPut_Key_3_756;
              verilogPut_Data_763 <= verilogPut_Data_3_759;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        956: begin
          if (verilogPut_index_768 == verilogPut_size_741) begin
            verilogPut_size_741 <= verilogPut_size_741+1;
          end
          case (verilogPut_index_768)
            0: begin
              verilogPut_Key_0_744 <= verilogPut_Key_761;
              verilogPut_Data_0_747 <= verilogPut_indexLeft_1473;
            end
            1: begin
              verilogPut_Key_1_748 <= verilogPut_Key_761;
              verilogPut_Data_1_751 <= verilogPut_indexLeft_1473;
            end
            2: begin
              verilogPut_Key_2_752 <= verilogPut_Key_761;
              verilogPut_Data_2_755 <= verilogPut_indexLeft_1473;
            end
            3: begin
              verilogPut_Key_3_756 <= verilogPut_Key_761;
              verilogPut_Data_3_759 <= verilogPut_indexLeft_1473;
            end
          endcase
          verilogPut_pc <= verilogPut_pc + 1;
        end
        957: begin
          verilogPut_success_1476 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        958: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_1415;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_1416;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_1415;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_1419;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_1423;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_1427;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_1431;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_1415;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_1422;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_1426;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_1430;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_1434;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        959: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        960: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        961: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        962: begin
          verilogPut_stuckSize_6_index_35 <= verilogPut_index_740;
          verilogPut_stuckSize_6_value_36 <= verilogPut_size_741;
          stuckSize_6_requestedAt <= step;
          verilogPut_stuckKeys_2_index_23 <= verilogPut_index_740;
          verilogPut_stuckKeys_2_value_24 <= verilogPut_Key_0_744;
          verilogPut_stuckKeys_2_value_25 <= verilogPut_Key_1_748;
          verilogPut_stuckKeys_2_value_26 <= verilogPut_Key_2_752;
          verilogPut_stuckKeys_2_value_27 <= verilogPut_Key_3_756;
          stuckKeys_2_requestedAt <= step;
          verilogPut_stuckData_4_index_29 <= verilogPut_index_740;
          verilogPut_stuckData_4_value_30 <= verilogPut_Data_0_747;
          verilogPut_stuckData_4_value_31 <= verilogPut_Data_1_751;
          verilogPut_stuckData_4_value_32 <= verilogPut_Data_2_755;
          verilogPut_stuckData_4_value_33 <= verilogPut_Data_3_759;
          stuckData_4_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        963: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        964: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        965: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        966: begin
          verilogPut_root_1479 <= 0;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        967: begin
          verilogPut_freeNext_9_index_192 <= verilogPut_root_1479;
          freeNext_9_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        968: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        969: begin
          verilogPut_next_1478 <= freeNext_freeNext_9_result_0;
          verilogPut_freeNext_10_index_193 <= verilogPut_root_1479;
          verilogPut_freeNext_10_value_194 <= verilogPut_indexRight_1474;
          freeNext_10_requestedAt <= step;
          verilogPut_isFree_1480 <= 1;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        970: begin
          verilogPut_stuckIsFree_11_index_195 <= verilogPut_indexRight_1474;
          verilogPut_stuckIsFree_11_value_196 <= verilogPut_isFree_1480;
          stuckIsFree_11_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        971: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        972: begin
          verilogPut_freeNext_10_index_193 <= verilogPut_indexRight_1474;
          verilogPut_freeNext_10_value_194 <= verilogPut_next_1478;
          freeNext_10_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        973: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        974: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        975: begin
          verilogPut_pc <= 976;
        end
        976: begin
          verilogPut_pc <= 977;
        end
        977: begin
          verilogPut_index_740 <= verilogPut_position_767;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        978: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        979: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        980: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        981: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        982: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        983: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        984: begin
          verilogPut_KeyCompares_0_745 <= verilogPut_k_0 <= verilogPut_Key_0_744 && 0 < verilogPut_size_741;
          verilogPut_KeyCollapse_0_746 <= 0;
          verilogPut_KeyCompares_1_749 <= verilogPut_k_0 >  verilogPut_Key_0_744 && verilogPut_k_0 <= verilogPut_Key_1_748 && 1 < verilogPut_size_741;
          verilogPut_KeyCollapse_1_750 <= 1;
          verilogPut_KeyCompares_2_753 <= verilogPut_k_0 >  verilogPut_Key_1_748 && verilogPut_k_0 <= verilogPut_Key_2_752 && 2 < verilogPut_size_741;
          verilogPut_KeyCollapse_2_754 <= 2;
          verilogPut_KeyCompares_3_757 <= verilogPut_k_0 >  verilogPut_Key_2_752 && verilogPut_k_0 <= verilogPut_Key_3_756 && 3 < verilogPut_size_741;
          verilogPut_KeyCollapse_3_758 <= 3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        985: begin
          if (verilogPut_KeyCompares_1_749) begin
            verilogPut_KeyCompares_0_745 <= 1;
            verilogPut_KeyCollapse_0_746 <= verilogPut_KeyCollapse_1_750;
          end
          if (verilogPut_KeyCompares_3_757) begin
            verilogPut_KeyCompares_2_753 <= 1;
            verilogPut_KeyCollapse_2_754 <= verilogPut_KeyCollapse_3_758;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        986: begin
          if (verilogPut_KeyCompares_2_753) begin
            verilogPut_KeyCompares_0_745 <= 1;
            verilogPut_KeyCollapse_0_746 <= verilogPut_KeyCollapse_2_754;
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        987: begin
          if (verilogPut_KeyCompares_0_745) begin
            verilogPut_Found_760 <= 1;
            case (verilogPut_KeyCollapse_0_746)
              0: begin
                verilogPut_StuckIndex_765 <= 0;
                verilogPut_FoundKey_762 <= verilogPut_Key_0_744;
                verilogPut_Data_763 <= verilogPut_Data_0_747;
              end
              1: begin
                verilogPut_StuckIndex_765 <= 1;
                verilogPut_FoundKey_762 <= verilogPut_Key_1_748;
                verilogPut_Data_763 <= verilogPut_Data_1_751;
              end
              2: begin
                verilogPut_StuckIndex_765 <= 2;
                verilogPut_FoundKey_762 <= verilogPut_Key_2_752;
                verilogPut_Data_763 <= verilogPut_Data_2_755;
              end
              3: begin
                verilogPut_StuckIndex_765 <= 3;
                verilogPut_FoundKey_762 <= verilogPut_Key_3_756;
                verilogPut_Data_763 <= verilogPut_Data_3_759;
              end
            endcase
          end
          else begin
            verilogPut_Found_760 <= 0;
            case (verilogPut_size_741)
              0: begin
                verilogPut_StuckIndex_765 <= 0;
                verilogPut_Data_763 <= verilogPut_Data_0_747;
              end
              1: begin
                verilogPut_StuckIndex_765 <= 1;
                verilogPut_Data_763 <= verilogPut_Data_1_751;
              end
              2: begin
                verilogPut_StuckIndex_765 <= 2;
                verilogPut_Data_763 <= verilogPut_Data_2_755;
              end
              3: begin
                verilogPut_StuckIndex_765 <= 3;
                verilogPut_Data_763 <= verilogPut_Data_3_759;
              end
            endcase
          end
          verilogPut_pc <= verilogPut_pc + 1;
        end
        988: begin
          verilogPut_position_767 <= verilogPut_Data_763;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        989: begin
          verilogPut_index_740 <= verilogPut_position_767;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        990: begin
          verilogPut_stuckSize_5_index_34 <= verilogPut_index_740;
          stuckSize_5_requestedAt <= step;
          verilogPut_stuckIsLeaf_7_index_37 <= verilogPut_index_740;
          stuckIsLeaf_7_requestedAt <= step;
          verilogPut_stuckKeys_1_index_22 <= verilogPut_index_740;
          stuckKeys_1_requestedAt <= step;
          verilogPut_stuckData_3_index_28 <= verilogPut_index_740;
          stuckData_3_requestedAt <= step;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        991: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        992: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        993: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        994: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        995: begin
          verilogPut_size_741 <= stuckSize_stuckSize_5_result_0;
          verilogPut_isLeaf_742 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          verilogPut_Key_0_744 <= stuckKeys_stuckKeys_1_result_0;
          verilogPut_Data_0_747 <= stuckData_stuckData_3_result_0;
          verilogPut_Key_1_748 <= stuckKeys_stuckKeys_1_result_1;
          verilogPut_Data_1_751 <= stuckData_stuckData_3_result_1;
          verilogPut_Key_2_752 <= stuckKeys_stuckKeys_1_result_2;
          verilogPut_Data_2_755 <= stuckData_stuckData_3_result_2;
          verilogPut_Key_3_756 <= stuckKeys_stuckKeys_1_result_3;
          verilogPut_Data_3_759 <= stuckData_stuckData_3_result_3;
          verilogPut_pc <= verilogPut_pc + 1;
        end
        996: begin
          if (verilogPut_isLeaf_742 == 0) begin
            verilogPut_pc <= 999;
          end
          else begin
            verilogPut_pc <= verilogPut_pc + 1;
          end
        end
        997: begin
          verilogPut_pc <= 1000;
        end
        998: begin
          verilogPut_pc <= 1000;
        end
        999: begin
          verilogPut_pc <= 586;
        end
        default: verilogPut_stop <= 1;
      endcase
    end
  end
endmodule
