//-----------------------------------------------------------------------------
// Database on a chip test bench
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree;                                                                      // Test bench for database on a chip
  reg                    stop;                                                  // Program has stopped when this goes high
  reg                   clock;                                                  // Clock
  integer                step;                                                  // Step of the simulation
  integer            maxSteps;                                                  // Maximum number of steps to execute
  integer          returnCode;                                                  // Return code
  integer      processCurrent;                                                  // To ensure we get the same results in Java and Verilog we have to run the processes single threaded in a constant order

  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_stop||stuckData_stop||put_stop;                                                             // Or of process stop fields

  initial begin
    returnCode = 0;
    maxSteps = 40000;
    for(step = -1; step < 0 || step < maxSteps && !stop; step = step + 1) begin // Steps below zero are run unconditionally to initialize each process so that Java and Verilog start in sync at step zero

      processCurrent = 0; clock = 0; #1; clock = 1; #1; // process_stuckIsLeaf_0000
      processCurrent = 1; clock = 0; #1; clock = 1; #1; // process_stuckIsFree_0001
      processCurrent = 2; clock = 0; #1; clock = 1; #1; // process_freeNext_0002
      processCurrent = 3; clock = 0; #1; clock = 1; #1; // process_stuckSize_0003
      processCurrent = 4; clock = 0; #1; clock = 1; #1; // process_stuckKeys_0004
      processCurrent = 5; clock = 0; #1; clock = 1; #1; // process_stuckData_0005
      processCurrent = 6; clock = 0; #1; clock = 1; #1; // process_put_0006
      if (step >= 0) chipPrint();                                            // Steps prior to zero are for initialization to make Java and Verilog match
    end
    if (!stop) $finish(1); else $finish(0);                                // Set return code depending on whether the simulation halted
  end
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[32*1];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_7_result_0;
  integer stuckIsLeaf_7_requestedAt;
  integer stuckIsLeaf_7_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_7_returnCode;
  integer stuckIsLeaf_8_requestedAt;
  integer stuckIsLeaf_8_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_8_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_7_result_0 <= 0;
      stuckIsLeaf_7_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_7_returnCode <= 0;
      stuckIsLeaf_8_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_8_returnCode <= 0;
      stuckIsLeaf_memory[0] <= 1;
      stuckIsLeaf_memory[1] <= 0;
      stuckIsLeaf_memory[2] <= 0;
      stuckIsLeaf_memory[3] <= 0;
      stuckIsLeaf_memory[4] <= 0;
      stuckIsLeaf_memory[5] <= 0;
      stuckIsLeaf_memory[6] <= 0;
      stuckIsLeaf_memory[7] <= 0;
      stuckIsLeaf_memory[8] <= 0;
      stuckIsLeaf_memory[9] <= 0;
      stuckIsLeaf_memory[10] <= 0;
      stuckIsLeaf_memory[11] <= 0;
      stuckIsLeaf_memory[12] <= 0;
      stuckIsLeaf_memory[13] <= 0;
      stuckIsLeaf_memory[14] <= 0;
      stuckIsLeaf_memory[15] <= 0;
      stuckIsLeaf_memory[16] <= 0;
      stuckIsLeaf_memory[17] <= 0;
      stuckIsLeaf_memory[18] <= 0;
      stuckIsLeaf_memory[19] <= 0;
      stuckIsLeaf_memory[20] <= 0;
      stuckIsLeaf_memory[21] <= 0;
      stuckIsLeaf_memory[22] <= 0;
      stuckIsLeaf_memory[23] <= 0;
      stuckIsLeaf_memory[24] <= 0;
      stuckIsLeaf_memory[25] <= 0;
      stuckIsLeaf_memory[26] <= 0;
      stuckIsLeaf_memory[27] <= 0;
      stuckIsLeaf_memory[28] <= 0;
      stuckIsLeaf_memory[29] <= 0;
      stuckIsLeaf_memory[30] <= 0;
      stuckIsLeaf_memory[31] <= 0;
    end
    else if (processCurrent == 0) begin
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_7_result_0 <= stuckIsLeaf_memory[put_stuckIsLeaf_7_index_39*1+0];
            stuckIsLeaf_7_finishedAt <= step;
          end
          else if ((stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step)) begin
            stuckIsLeaf_memory[put_stuckIsLeaf_8_index_40*1+0] <= put_stuckIsLeaf_8_value_41;
            stuckIsLeaf_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[32*1];
  integer stuckIsFree_11_requestedAt;
  integer stuckIsFree_11_finishedAt;
  integer stuckIsFree_stuckIsFree_11_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_11_finishedAt <= -1;
      stuckIsFree_stuckIsFree_11_returnCode <= 0;
      stuckIsFree_memory[0] <= 0;
      stuckIsFree_memory[1] <= 1;
      stuckIsFree_memory[2] <= 1;
      stuckIsFree_memory[3] <= 1;
      stuckIsFree_memory[4] <= 1;
      stuckIsFree_memory[5] <= 1;
      stuckIsFree_memory[6] <= 1;
      stuckIsFree_memory[7] <= 1;
      stuckIsFree_memory[8] <= 1;
      stuckIsFree_memory[9] <= 1;
      stuckIsFree_memory[10] <= 1;
      stuckIsFree_memory[11] <= 1;
      stuckIsFree_memory[12] <= 1;
      stuckIsFree_memory[13] <= 1;
      stuckIsFree_memory[14] <= 1;
      stuckIsFree_memory[15] <= 1;
      stuckIsFree_memory[16] <= 1;
      stuckIsFree_memory[17] <= 1;
      stuckIsFree_memory[18] <= 1;
      stuckIsFree_memory[19] <= 1;
      stuckIsFree_memory[20] <= 1;
      stuckIsFree_memory[21] <= 1;
      stuckIsFree_memory[22] <= 1;
      stuckIsFree_memory[23] <= 1;
      stuckIsFree_memory[24] <= 1;
      stuckIsFree_memory[25] <= 1;
      stuckIsFree_memory[26] <= 1;
      stuckIsFree_memory[27] <= 1;
      stuckIsFree_memory[28] <= 1;
      stuckIsFree_memory[29] <= 1;
      stuckIsFree_memory[30] <= 1;
      stuckIsFree_memory[31] <= 1;
    end
    else if (processCurrent == 1) begin
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step)) begin
            stuckIsFree_memory[put_stuckIsFree_11_index_197*1+0] <= put_stuckIsFree_11_value_198;
            stuckIsFree_11_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [6-1:0] freeNext_memory[32*1];
  reg [6-1:0] freeNext_freeNext_9_result_0;
  integer freeNext_9_requestedAt;
  integer freeNext_9_finishedAt;
  integer freeNext_freeNext_9_returnCode;
  integer freeNext_10_requestedAt;
  integer freeNext_10_finishedAt;
  integer freeNext_freeNext_10_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_9_result_0 <= 0;
      freeNext_9_finishedAt <= -1;
      freeNext_freeNext_9_returnCode <= 0;
      freeNext_10_finishedAt <= -1;
      freeNext_freeNext_10_returnCode <= 0;
      freeNext_memory[0] <= 1;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 7;
      freeNext_memory[7] <= 8;
      freeNext_memory[8] <= 9;
      freeNext_memory[9] <= 10;
      freeNext_memory[10] <= 11;
      freeNext_memory[11] <= 12;
      freeNext_memory[12] <= 13;
      freeNext_memory[13] <= 14;
      freeNext_memory[14] <= 15;
      freeNext_memory[15] <= 16;
      freeNext_memory[16] <= 17;
      freeNext_memory[17] <= 18;
      freeNext_memory[18] <= 19;
      freeNext_memory[19] <= 20;
      freeNext_memory[20] <= 21;
      freeNext_memory[21] <= 22;
      freeNext_memory[22] <= 23;
      freeNext_memory[23] <= 24;
      freeNext_memory[24] <= 25;
      freeNext_memory[25] <= 26;
      freeNext_memory[26] <= 27;
      freeNext_memory[27] <= 28;
      freeNext_memory[28] <= 29;
      freeNext_memory[29] <= 30;
      freeNext_memory[30] <= 31;
      freeNext_memory[31] <= 0;
    end
    else if (processCurrent == 2) begin
      case(freeNext_pc)
        0: begin
          if ((freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step)) begin
            freeNext_freeNext_9_result_0 <= freeNext_memory[put_freeNext_9_index_194*1+0];
            freeNext_9_finishedAt <= step;
          end
          else if ((freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step)) begin
            freeNext_memory[put_freeNext_10_index_195*1+0] <= put_freeNext_10_value_196;
            freeNext_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[32*1];
  reg [3-1:0] stuckSize_stuckSize_5_result_0;
  integer stuckSize_5_requestedAt;
  integer stuckSize_5_finishedAt;
  integer stuckSize_stuckSize_5_returnCode;
  integer stuckSize_6_requestedAt;
  integer stuckSize_6_finishedAt;
  integer stuckSize_stuckSize_6_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_5_result_0 <= 0;
      stuckSize_5_finishedAt <= -1;
      stuckSize_stuckSize_5_returnCode <= 0;
      stuckSize_6_finishedAt <= -1;
      stuckSize_stuckSize_6_returnCode <= 0;
      stuckSize_memory[0] <= 0;
      stuckSize_memory[1] <= 0;
      stuckSize_memory[2] <= 0;
      stuckSize_memory[3] <= 0;
      stuckSize_memory[4] <= 0;
      stuckSize_memory[5] <= 0;
      stuckSize_memory[6] <= 0;
      stuckSize_memory[7] <= 0;
      stuckSize_memory[8] <= 0;
      stuckSize_memory[9] <= 0;
      stuckSize_memory[10] <= 0;
      stuckSize_memory[11] <= 0;
      stuckSize_memory[12] <= 0;
      stuckSize_memory[13] <= 0;
      stuckSize_memory[14] <= 0;
      stuckSize_memory[15] <= 0;
      stuckSize_memory[16] <= 0;
      stuckSize_memory[17] <= 0;
      stuckSize_memory[18] <= 0;
      stuckSize_memory[19] <= 0;
      stuckSize_memory[20] <= 0;
      stuckSize_memory[21] <= 0;
      stuckSize_memory[22] <= 0;
      stuckSize_memory[23] <= 0;
      stuckSize_memory[24] <= 0;
      stuckSize_memory[25] <= 0;
      stuckSize_memory[26] <= 0;
      stuckSize_memory[27] <= 0;
      stuckSize_memory[28] <= 0;
      stuckSize_memory[29] <= 0;
      stuckSize_memory[30] <= 0;
      stuckSize_memory[31] <= 0;
    end
    else if (processCurrent == 3) begin
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step)) begin
            stuckSize_stuckSize_5_result_0 <= stuckSize_memory[put_stuckSize_5_index_36*1+0];
            stuckSize_5_finishedAt <= step;
          end
          else if ((stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step)) begin
            stuckSize_memory[put_stuckSize_6_index_37*1+0] <= put_stuckSize_6_value_38;
            stuckSize_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys  process_stuckKeys_0004
  (* ram_style = "block" *)
  reg [8-1:0] stuckKeys_memory[32*4];
  reg [8-1:0] stuckKeys_stuckKeys_1_result_0;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_1;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_2;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_3;
  integer stuckKeys_1_requestedAt;
  integer stuckKeys_1_finishedAt;
  integer stuckKeys_stuckKeys_1_returnCode;
  integer stuckKeys_2_requestedAt;
  integer stuckKeys_2_finishedAt;
  integer stuckKeys_stuckKeys_2_returnCode;
  integer stuckKeys_pc;
  integer stuckKeys_stop;
  integer stuckKeys_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_pc <= 0;
      stuckKeys_stop <= 0;
      stuckKeys_returnCode <= 0;
      stuckKeys_stuckKeys_1_result_0 <= 0;
      stuckKeys_stuckKeys_1_result_1 <= 0;
      stuckKeys_stuckKeys_1_result_2 <= 0;
      stuckKeys_stuckKeys_1_result_3 <= 0;
      stuckKeys_1_finishedAt <= -1;
      stuckKeys_stuckKeys_1_returnCode <= 0;
      stuckKeys_2_finishedAt <= -1;
      stuckKeys_stuckKeys_2_returnCode <= 0;
      stuckKeys_memory[0] <= 0;
      stuckKeys_memory[1] <= 0;
      stuckKeys_memory[2] <= 0;
      stuckKeys_memory[3] <= 0;
      stuckKeys_memory[4] <= 0;
      stuckKeys_memory[5] <= 0;
      stuckKeys_memory[6] <= 0;
      stuckKeys_memory[7] <= 0;
      stuckKeys_memory[8] <= 0;
      stuckKeys_memory[9] <= 0;
      stuckKeys_memory[10] <= 0;
      stuckKeys_memory[11] <= 0;
      stuckKeys_memory[12] <= 0;
      stuckKeys_memory[13] <= 0;
      stuckKeys_memory[14] <= 0;
      stuckKeys_memory[15] <= 0;
      stuckKeys_memory[16] <= 0;
      stuckKeys_memory[17] <= 0;
      stuckKeys_memory[18] <= 0;
      stuckKeys_memory[19] <= 0;
      stuckKeys_memory[20] <= 0;
      stuckKeys_memory[21] <= 0;
      stuckKeys_memory[22] <= 0;
      stuckKeys_memory[23] <= 0;
      stuckKeys_memory[24] <= 0;
      stuckKeys_memory[25] <= 0;
      stuckKeys_memory[26] <= 0;
      stuckKeys_memory[27] <= 0;
      stuckKeys_memory[28] <= 0;
      stuckKeys_memory[29] <= 0;
      stuckKeys_memory[30] <= 0;
      stuckKeys_memory[31] <= 0;
      stuckKeys_memory[32] <= 0;
      stuckKeys_memory[33] <= 0;
      stuckKeys_memory[34] <= 0;
      stuckKeys_memory[35] <= 0;
      stuckKeys_memory[36] <= 0;
      stuckKeys_memory[37] <= 0;
      stuckKeys_memory[38] <= 0;
      stuckKeys_memory[39] <= 0;
      stuckKeys_memory[40] <= 0;
      stuckKeys_memory[41] <= 0;
      stuckKeys_memory[42] <= 0;
      stuckKeys_memory[43] <= 0;
      stuckKeys_memory[44] <= 0;
      stuckKeys_memory[45] <= 0;
      stuckKeys_memory[46] <= 0;
      stuckKeys_memory[47] <= 0;
      stuckKeys_memory[48] <= 0;
      stuckKeys_memory[49] <= 0;
      stuckKeys_memory[50] <= 0;
      stuckKeys_memory[51] <= 0;
      stuckKeys_memory[52] <= 0;
      stuckKeys_memory[53] <= 0;
      stuckKeys_memory[54] <= 0;
      stuckKeys_memory[55] <= 0;
      stuckKeys_memory[56] <= 0;
      stuckKeys_memory[57] <= 0;
      stuckKeys_memory[58] <= 0;
      stuckKeys_memory[59] <= 0;
      stuckKeys_memory[60] <= 0;
      stuckKeys_memory[61] <= 0;
      stuckKeys_memory[62] <= 0;
      stuckKeys_memory[63] <= 0;
      stuckKeys_memory[64] <= 0;
      stuckKeys_memory[65] <= 0;
      stuckKeys_memory[66] <= 0;
      stuckKeys_memory[67] <= 0;
      stuckKeys_memory[68] <= 0;
      stuckKeys_memory[69] <= 0;
      stuckKeys_memory[70] <= 0;
      stuckKeys_memory[71] <= 0;
      stuckKeys_memory[72] <= 0;
      stuckKeys_memory[73] <= 0;
      stuckKeys_memory[74] <= 0;
      stuckKeys_memory[75] <= 0;
      stuckKeys_memory[76] <= 0;
      stuckKeys_memory[77] <= 0;
      stuckKeys_memory[78] <= 0;
      stuckKeys_memory[79] <= 0;
      stuckKeys_memory[80] <= 0;
      stuckKeys_memory[81] <= 0;
      stuckKeys_memory[82] <= 0;
      stuckKeys_memory[83] <= 0;
      stuckKeys_memory[84] <= 0;
      stuckKeys_memory[85] <= 0;
      stuckKeys_memory[86] <= 0;
      stuckKeys_memory[87] <= 0;
      stuckKeys_memory[88] <= 0;
      stuckKeys_memory[89] <= 0;
      stuckKeys_memory[90] <= 0;
      stuckKeys_memory[91] <= 0;
      stuckKeys_memory[92] <= 0;
      stuckKeys_memory[93] <= 0;
      stuckKeys_memory[94] <= 0;
      stuckKeys_memory[95] <= 0;
      stuckKeys_memory[96] <= 0;
      stuckKeys_memory[97] <= 0;
      stuckKeys_memory[98] <= 0;
      stuckKeys_memory[99] <= 0;
      stuckKeys_memory[100] <= 0;
      stuckKeys_memory[101] <= 0;
      stuckKeys_memory[102] <= 0;
      stuckKeys_memory[103] <= 0;
      stuckKeys_memory[104] <= 0;
      stuckKeys_memory[105] <= 0;
      stuckKeys_memory[106] <= 0;
      stuckKeys_memory[107] <= 0;
      stuckKeys_memory[108] <= 0;
      stuckKeys_memory[109] <= 0;
      stuckKeys_memory[110] <= 0;
      stuckKeys_memory[111] <= 0;
      stuckKeys_memory[112] <= 0;
      stuckKeys_memory[113] <= 0;
      stuckKeys_memory[114] <= 0;
      stuckKeys_memory[115] <= 0;
      stuckKeys_memory[116] <= 0;
      stuckKeys_memory[117] <= 0;
      stuckKeys_memory[118] <= 0;
      stuckKeys_memory[119] <= 0;
      stuckKeys_memory[120] <= 0;
      stuckKeys_memory[121] <= 0;
      stuckKeys_memory[122] <= 0;
      stuckKeys_memory[123] <= 0;
      stuckKeys_memory[124] <= 0;
      stuckKeys_memory[125] <= 0;
      stuckKeys_memory[126] <= 0;
      stuckKeys_memory[127] <= 0;
    end
    else if (processCurrent == 4) begin
      case(stuckKeys_pc)
        0: begin
          if ((stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step)) begin
            stuckKeys_stuckKeys_1_result_0 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+0];
            stuckKeys_stuckKeys_1_result_1 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+1];
            stuckKeys_stuckKeys_1_result_2 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+2];
            stuckKeys_stuckKeys_1_result_3 <= stuckKeys_memory[put_stuckKeys_1_index_24*4+3];
            stuckKeys_1_finishedAt <= step;
          end
          else if ((stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step)) begin
            stuckKeys_memory[put_stuckKeys_2_index_25*4+0] <= put_stuckKeys_2_value_26;
            stuckKeys_memory[put_stuckKeys_2_index_25*4+1] <= put_stuckKeys_2_value_27;
            stuckKeys_memory[put_stuckKeys_2_index_25*4+2] <= put_stuckKeys_2_value_28;
            stuckKeys_memory[put_stuckKeys_2_index_25*4+3] <= put_stuckKeys_2_value_29;
            stuckKeys_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_stop <= 1;
      endcase
    end
  end
  // Process: stuckData  process_stuckData_0005
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_memory[32*4];
  reg [8-1:0] stuckData_stuckData_3_result_0;
  reg [8-1:0] stuckData_stuckData_3_result_1;
  reg [8-1:0] stuckData_stuckData_3_result_2;
  reg [8-1:0] stuckData_stuckData_3_result_3;
  integer stuckData_3_requestedAt;
  integer stuckData_3_finishedAt;
  integer stuckData_stuckData_3_returnCode;
  integer stuckData_4_requestedAt;
  integer stuckData_4_finishedAt;
  integer stuckData_stuckData_4_returnCode;
  integer stuckData_pc;
  integer stuckData_stop;
  integer stuckData_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_pc <= 0;
      stuckData_stop <= 0;
      stuckData_returnCode <= 0;
      stuckData_stuckData_3_result_0 <= 0;
      stuckData_stuckData_3_result_1 <= 0;
      stuckData_stuckData_3_result_2 <= 0;
      stuckData_stuckData_3_result_3 <= 0;
      stuckData_3_finishedAt <= -1;
      stuckData_stuckData_3_returnCode <= 0;
      stuckData_4_finishedAt <= -1;
      stuckData_stuckData_4_returnCode <= 0;
      stuckData_memory[0] <= 0;
      stuckData_memory[1] <= 0;
      stuckData_memory[2] <= 0;
      stuckData_memory[3] <= 0;
      stuckData_memory[4] <= 0;
      stuckData_memory[5] <= 0;
      stuckData_memory[6] <= 0;
      stuckData_memory[7] <= 0;
      stuckData_memory[8] <= 0;
      stuckData_memory[9] <= 0;
      stuckData_memory[10] <= 0;
      stuckData_memory[11] <= 0;
      stuckData_memory[12] <= 0;
      stuckData_memory[13] <= 0;
      stuckData_memory[14] <= 0;
      stuckData_memory[15] <= 0;
      stuckData_memory[16] <= 0;
      stuckData_memory[17] <= 0;
      stuckData_memory[18] <= 0;
      stuckData_memory[19] <= 0;
      stuckData_memory[20] <= 0;
      stuckData_memory[21] <= 0;
      stuckData_memory[22] <= 0;
      stuckData_memory[23] <= 0;
      stuckData_memory[24] <= 0;
      stuckData_memory[25] <= 0;
      stuckData_memory[26] <= 0;
      stuckData_memory[27] <= 0;
      stuckData_memory[28] <= 0;
      stuckData_memory[29] <= 0;
      stuckData_memory[30] <= 0;
      stuckData_memory[31] <= 0;
      stuckData_memory[32] <= 0;
      stuckData_memory[33] <= 0;
      stuckData_memory[34] <= 0;
      stuckData_memory[35] <= 0;
      stuckData_memory[36] <= 0;
      stuckData_memory[37] <= 0;
      stuckData_memory[38] <= 0;
      stuckData_memory[39] <= 0;
      stuckData_memory[40] <= 0;
      stuckData_memory[41] <= 0;
      stuckData_memory[42] <= 0;
      stuckData_memory[43] <= 0;
      stuckData_memory[44] <= 0;
      stuckData_memory[45] <= 0;
      stuckData_memory[46] <= 0;
      stuckData_memory[47] <= 0;
      stuckData_memory[48] <= 0;
      stuckData_memory[49] <= 0;
      stuckData_memory[50] <= 0;
      stuckData_memory[51] <= 0;
      stuckData_memory[52] <= 0;
      stuckData_memory[53] <= 0;
      stuckData_memory[54] <= 0;
      stuckData_memory[55] <= 0;
      stuckData_memory[56] <= 0;
      stuckData_memory[57] <= 0;
      stuckData_memory[58] <= 0;
      stuckData_memory[59] <= 0;
      stuckData_memory[60] <= 0;
      stuckData_memory[61] <= 0;
      stuckData_memory[62] <= 0;
      stuckData_memory[63] <= 0;
      stuckData_memory[64] <= 0;
      stuckData_memory[65] <= 0;
      stuckData_memory[66] <= 0;
      stuckData_memory[67] <= 0;
      stuckData_memory[68] <= 0;
      stuckData_memory[69] <= 0;
      stuckData_memory[70] <= 0;
      stuckData_memory[71] <= 0;
      stuckData_memory[72] <= 0;
      stuckData_memory[73] <= 0;
      stuckData_memory[74] <= 0;
      stuckData_memory[75] <= 0;
      stuckData_memory[76] <= 0;
      stuckData_memory[77] <= 0;
      stuckData_memory[78] <= 0;
      stuckData_memory[79] <= 0;
      stuckData_memory[80] <= 0;
      stuckData_memory[81] <= 0;
      stuckData_memory[82] <= 0;
      stuckData_memory[83] <= 0;
      stuckData_memory[84] <= 0;
      stuckData_memory[85] <= 0;
      stuckData_memory[86] <= 0;
      stuckData_memory[87] <= 0;
      stuckData_memory[88] <= 0;
      stuckData_memory[89] <= 0;
      stuckData_memory[90] <= 0;
      stuckData_memory[91] <= 0;
      stuckData_memory[92] <= 0;
      stuckData_memory[93] <= 0;
      stuckData_memory[94] <= 0;
      stuckData_memory[95] <= 0;
      stuckData_memory[96] <= 0;
      stuckData_memory[97] <= 0;
      stuckData_memory[98] <= 0;
      stuckData_memory[99] <= 0;
      stuckData_memory[100] <= 0;
      stuckData_memory[101] <= 0;
      stuckData_memory[102] <= 0;
      stuckData_memory[103] <= 0;
      stuckData_memory[104] <= 0;
      stuckData_memory[105] <= 0;
      stuckData_memory[106] <= 0;
      stuckData_memory[107] <= 0;
      stuckData_memory[108] <= 0;
      stuckData_memory[109] <= 0;
      stuckData_memory[110] <= 0;
      stuckData_memory[111] <= 0;
      stuckData_memory[112] <= 0;
      stuckData_memory[113] <= 0;
      stuckData_memory[114] <= 0;
      stuckData_memory[115] <= 0;
      stuckData_memory[116] <= 0;
      stuckData_memory[117] <= 0;
      stuckData_memory[118] <= 0;
      stuckData_memory[119] <= 0;
      stuckData_memory[120] <= 0;
      stuckData_memory[121] <= 0;
      stuckData_memory[122] <= 0;
      stuckData_memory[123] <= 0;
      stuckData_memory[124] <= 0;
      stuckData_memory[125] <= 0;
      stuckData_memory[126] <= 0;
      stuckData_memory[127] <= 0;
    end
    else if (processCurrent == 5) begin
      case(stuckData_pc)
        0: begin
          if ((stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step)) begin
            stuckData_stuckData_3_result_0 <= stuckData_memory[put_stuckData_3_index_30*4+0];
            stuckData_stuckData_3_result_1 <= stuckData_memory[put_stuckData_3_index_30*4+1];
            stuckData_stuckData_3_result_2 <= stuckData_memory[put_stuckData_3_index_30*4+2];
            stuckData_stuckData_3_result_3 <= stuckData_memory[put_stuckData_3_index_30*4+3];
            stuckData_3_finishedAt <= step;
          end
          else if ((stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step)) begin
            stuckData_memory[put_stuckData_4_index_31*4+0] <= put_stuckData_4_value_32;
            stuckData_memory[put_stuckData_4_index_31*4+1] <= put_stuckData_4_value_33;
            stuckData_memory[put_stuckData_4_index_31*4+2] <= put_stuckData_4_value_34;
            stuckData_memory[put_stuckData_4_index_31*4+3] <= put_stuckData_4_value_35;
            stuckData_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_stop <= 1;
      endcase
    end
  end
  // Process: put  process_put_0006
  reg [8-1:0] put_k_0;
  reg [8-1:0] put_d_1;
  reg [8-1:0] put_i_2;
  reg [1-1:0] put_l_3;
  reg [6-1:0] put_index_4;
  reg [3-1:0] put_size_5;
  reg [1-1:0] put_isLeaf_6;
  reg [6-1:0] put_nextFree_7;
  reg [8-1:0] put_Key_0_8;
  reg [1-1:0] put_KeyCompares_0_9;
  reg [3-1:0] put_KeyCollapse_0_10;
  reg [8-1:0] put_Data_0_11;
  reg [8-1:0] put_Key_1_12;
  reg [1-1:0] put_KeyCompares_1_13;
  reg [3-1:0] put_KeyCollapse_1_14;
  reg [8-1:0] put_Data_1_15;
  reg [8-1:0] put_Key_2_16;
  reg [1-1:0] put_KeyCompares_2_17;
  reg [3-1:0] put_KeyCollapse_2_18;
  reg [8-1:0] put_Data_2_19;
  reg [8-1:0] put_Key_3_20;
  reg [1-1:0] put_KeyCompares_3_21;
  reg [3-1:0] put_KeyCollapse_3_22;
  reg [8-1:0] put_Data_3_23;
  reg [5-1:0] put_stuckKeys_1_index_24;
  reg [5-1:0] put_stuckKeys_2_index_25;
  reg [8-1:0] put_stuckKeys_2_value_26;
  reg [8-1:0] put_stuckKeys_2_value_27;
  reg [8-1:0] put_stuckKeys_2_value_28;
  reg [8-1:0] put_stuckKeys_2_value_29;
  reg [5-1:0] put_stuckData_3_index_30;
  reg [5-1:0] put_stuckData_4_index_31;
  reg [8-1:0] put_stuckData_4_value_32;
  reg [8-1:0] put_stuckData_4_value_33;
  reg [8-1:0] put_stuckData_4_value_34;
  reg [8-1:0] put_stuckData_4_value_35;
  reg [5-1:0] put_stuckSize_5_index_36;
  reg [5-1:0] put_stuckSize_6_index_37;
  reg [3-1:0] put_stuckSize_6_value_38;
  reg [5-1:0] put_stuckIsLeaf_7_index_39;
  reg [5-1:0] put_stuckIsLeaf_8_index_40;
  reg [1-1:0] put_stuckIsLeaf_8_value_41;
  reg [1-1:0] put_Found_42;
  reg [8-1:0] put_Key_43;
  reg [8-1:0] put_FoundKey_44;
  reg [8-1:0] put_Data_45;
  reg [6-1:0] put_BtreeIndex_46;
  reg [3-1:0] put_StuckIndex_47;
  reg [1-1:0] put_MergeSuccess_48;
  reg [6-1:0] put_index_49;
  reg [3-1:0] put_size_50;
  reg [1-1:0] put_isLeaf_51;
  reg [6-1:0] put_nextFree_52;
  reg [8-1:0] put_Key_0_53;
  reg [1-1:0] put_KeyCompares_0_54;
  reg [3-1:0] put_KeyCollapse_0_55;
  reg [8-1:0] put_Data_0_56;
  reg [8-1:0] put_Key_1_57;
  reg [1-1:0] put_KeyCompares_1_58;
  reg [3-1:0] put_KeyCollapse_1_59;
  reg [8-1:0] put_Data_1_60;
  reg [8-1:0] put_Key_2_61;
  reg [1-1:0] put_KeyCompares_2_62;
  reg [3-1:0] put_KeyCollapse_2_63;
  reg [8-1:0] put_Data_2_64;
  reg [8-1:0] put_Key_3_65;
  reg [1-1:0] put_KeyCompares_3_66;
  reg [3-1:0] put_KeyCollapse_3_67;
  reg [8-1:0] put_Data_3_68;
  reg [1-1:0] put_Found_69;
  reg [8-1:0] put_Key_70;
  reg [8-1:0] put_FoundKey_71;
  reg [8-1:0] put_Data_72;
  reg [6-1:0] put_BtreeIndex_73;
  reg [3-1:0] put_StuckIndex_74;
  reg [1-1:0] put_MergeSuccess_75;
  reg [6-1:0] put_index_76;
  reg [3-1:0] put_size_77;
  reg [1-1:0] put_isLeaf_78;
  reg [6-1:0] put_nextFree_79;
  reg [8-1:0] put_Key_0_80;
  reg [1-1:0] put_KeyCompares_0_81;
  reg [3-1:0] put_KeyCollapse_0_82;
  reg [8-1:0] put_Data_0_83;
  reg [8-1:0] put_Key_1_84;
  reg [1-1:0] put_KeyCompares_1_85;
  reg [3-1:0] put_KeyCollapse_1_86;
  reg [8-1:0] put_Data_1_87;
  reg [8-1:0] put_Key_2_88;
  reg [1-1:0] put_KeyCompares_2_89;
  reg [3-1:0] put_KeyCollapse_2_90;
  reg [8-1:0] put_Data_2_91;
  reg [8-1:0] put_Key_3_92;
  reg [1-1:0] put_KeyCompares_3_93;
  reg [3-1:0] put_KeyCollapse_3_94;
  reg [8-1:0] put_Data_3_95;
  reg [1-1:0] put_Found_96;
  reg [8-1:0] put_Key_97;
  reg [8-1:0] put_FoundKey_98;
  reg [8-1:0] put_Data_99;
  reg [6-1:0] put_BtreeIndex_100;
  reg [3-1:0] put_StuckIndex_101;
  reg [1-1:0] put_MergeSuccess_102;
  reg [6-1:0] put_child_103;
  reg [6-1:0] put_parent_104;
  reg [3-1:0] put_childInparent_105;
  reg [1-1:0] put_found_106;
  reg [1-1:0] put_full_107;
  reg [3-1:0] put_i_108;
  reg [1-1:0] put_notFull_109;
  reg [6-1:0] put_index_110;
  reg [3-1:0] put_size_111;
  reg [1-1:0] put_isLeaf_112;
  reg [6-1:0] put_nextFree_113;
  reg [8-1:0] put_Key_0_114;
  reg [1-1:0] put_KeyCompares_0_115;
  reg [3-1:0] put_KeyCollapse_0_116;
  reg [8-1:0] put_Data_0_117;
  reg [8-1:0] put_Key_1_118;
  reg [1-1:0] put_KeyCompares_1_119;
  reg [3-1:0] put_KeyCollapse_1_120;
  reg [8-1:0] put_Data_1_121;
  reg [8-1:0] put_Key_2_122;
  reg [1-1:0] put_KeyCompares_2_123;
  reg [3-1:0] put_KeyCollapse_2_124;
  reg [8-1:0] put_Data_2_125;
  reg [8-1:0] put_Key_3_126;
  reg [1-1:0] put_KeyCompares_3_127;
  reg [3-1:0] put_KeyCollapse_3_128;
  reg [8-1:0] put_Data_3_129;
  reg [1-1:0] put_Found_130;
  reg [8-1:0] put_Key_131;
  reg [8-1:0] put_FoundKey_132;
  reg [8-1:0] put_Data_133;
  reg [6-1:0] put_BtreeIndex_134;
  reg [3-1:0] put_StuckIndex_135;
  reg [1-1:0] put_MergeSuccess_136;
  reg [6-1:0] put_index_137;
  reg [3-1:0] put_size_138;
  reg [1-1:0] put_isLeaf_139;
  reg [6-1:0] put_nextFree_140;
  reg [8-1:0] put_Key_0_141;
  reg [1-1:0] put_KeyCompares_0_142;
  reg [3-1:0] put_KeyCollapse_0_143;
  reg [8-1:0] put_Data_0_144;
  reg [8-1:0] put_Key_1_145;
  reg [1-1:0] put_KeyCompares_1_146;
  reg [3-1:0] put_KeyCollapse_1_147;
  reg [8-1:0] put_Data_1_148;
  reg [8-1:0] put_Key_2_149;
  reg [1-1:0] put_KeyCompares_2_150;
  reg [3-1:0] put_KeyCollapse_2_151;
  reg [8-1:0] put_Data_2_152;
  reg [8-1:0] put_Key_3_153;
  reg [1-1:0] put_KeyCompares_3_154;
  reg [3-1:0] put_KeyCollapse_3_155;
  reg [8-1:0] put_Data_3_156;
  reg [1-1:0] put_Found_157;
  reg [8-1:0] put_Key_158;
  reg [8-1:0] put_FoundKey_159;
  reg [8-1:0] put_Data_160;
  reg [6-1:0] put_BtreeIndex_161;
  reg [3-1:0] put_StuckIndex_162;
  reg [1-1:0] put_MergeSuccess_163;
  reg [6-1:0] put_index_164;
  reg [3-1:0] put_size_165;
  reg [1-1:0] put_isLeaf_166;
  reg [6-1:0] put_nextFree_167;
  reg [8-1:0] put_Key_0_168;
  reg [1-1:0] put_KeyCompares_0_169;
  reg [3-1:0] put_KeyCollapse_0_170;
  reg [8-1:0] put_Data_0_171;
  reg [8-1:0] put_Key_1_172;
  reg [1-1:0] put_KeyCompares_1_173;
  reg [3-1:0] put_KeyCollapse_1_174;
  reg [8-1:0] put_Data_1_175;
  reg [8-1:0] put_Key_2_176;
  reg [1-1:0] put_KeyCompares_2_177;
  reg [3-1:0] put_KeyCollapse_2_178;
  reg [8-1:0] put_Data_2_179;
  reg [8-1:0] put_Key_3_180;
  reg [1-1:0] put_KeyCompares_3_181;
  reg [3-1:0] put_KeyCollapse_3_182;
  reg [8-1:0] put_Data_3_183;
  reg [1-1:0] put_Found_184;
  reg [8-1:0] put_Key_185;
  reg [8-1:0] put_FoundKey_186;
  reg [8-1:0] put_Data_187;
  reg [6-1:0] put_BtreeIndex_188;
  reg [3-1:0] put_StuckIndex_189;
  reg [1-1:0] put_MergeSuccess_190;
  reg [6-1:0] put_indexLeft_191;
  reg [6-1:0] put_indexRight_192;
  reg [8-1:0] put_midKey_193;
  reg [5-1:0] put_freeNext_9_index_194;
  reg [5-1:0] put_freeNext_10_index_195;
  reg [6-1:0] put_freeNext_10_value_196;
  reg [5-1:0] put_stuckIsFree_11_index_197;
  reg [1-1:0] put_stuckIsFree_11_value_198;
  reg [6-1:0] put_root_199;
  reg [6-1:0] put_next_200;
  reg [1-1:0] put_isLeaf_201;
  reg [1-1:0] put_isFree_202;
  reg [6-1:0] put_root_203;
  reg [6-1:0] put_next_204;
  reg [1-1:0] put_isLeaf_205;
  reg [1-1:0] put_isFree_206;
  reg [3-1:0] put_i_207;
  reg [1-1:0] put_notFull_208;
  reg [6-1:0] put_index_209;
  reg [3-1:0] put_size_210;
  reg [1-1:0] put_isLeaf_211;
  reg [6-1:0] put_nextFree_212;
  reg [8-1:0] put_Key_0_213;
  reg [1-1:0] put_KeyCompares_0_214;
  reg [3-1:0] put_KeyCollapse_0_215;
  reg [8-1:0] put_Data_0_216;
  reg [8-1:0] put_Key_1_217;
  reg [1-1:0] put_KeyCompares_1_218;
  reg [3-1:0] put_KeyCollapse_1_219;
  reg [8-1:0] put_Data_1_220;
  reg [8-1:0] put_Key_2_221;
  reg [1-1:0] put_KeyCompares_2_222;
  reg [3-1:0] put_KeyCollapse_2_223;
  reg [8-1:0] put_Data_2_224;
  reg [8-1:0] put_Key_3_225;
  reg [1-1:0] put_KeyCompares_3_226;
  reg [3-1:0] put_KeyCollapse_3_227;
  reg [8-1:0] put_Data_3_228;
  reg [1-1:0] put_Found_229;
  reg [8-1:0] put_Key_230;
  reg [8-1:0] put_FoundKey_231;
  reg [8-1:0] put_Data_232;
  reg [6-1:0] put_BtreeIndex_233;
  reg [3-1:0] put_StuckIndex_234;
  reg [1-1:0] put_MergeSuccess_235;
  reg [6-1:0] put_index_236;
  reg [3-1:0] put_size_237;
  reg [1-1:0] put_isLeaf_238;
  reg [6-1:0] put_nextFree_239;
  reg [8-1:0] put_Key_0_240;
  reg [1-1:0] put_KeyCompares_0_241;
  reg [3-1:0] put_KeyCollapse_0_242;
  reg [8-1:0] put_Data_0_243;
  reg [8-1:0] put_Key_1_244;
  reg [1-1:0] put_KeyCompares_1_245;
  reg [3-1:0] put_KeyCollapse_1_246;
  reg [8-1:0] put_Data_1_247;
  reg [8-1:0] put_Key_2_248;
  reg [1-1:0] put_KeyCompares_2_249;
  reg [3-1:0] put_KeyCollapse_2_250;
  reg [8-1:0] put_Data_2_251;
  reg [8-1:0] put_Key_3_252;
  reg [1-1:0] put_KeyCompares_3_253;
  reg [3-1:0] put_KeyCollapse_3_254;
  reg [8-1:0] put_Data_3_255;
  reg [1-1:0] put_Found_256;
  reg [8-1:0] put_Key_257;
  reg [8-1:0] put_FoundKey_258;
  reg [8-1:0] put_Data_259;
  reg [6-1:0] put_BtreeIndex_260;
  reg [3-1:0] put_StuckIndex_261;
  reg [1-1:0] put_MergeSuccess_262;
  reg [6-1:0] put_index_263;
  reg [3-1:0] put_size_264;
  reg [1-1:0] put_isLeaf_265;
  reg [6-1:0] put_nextFree_266;
  reg [8-1:0] put_Key_0_267;
  reg [1-1:0] put_KeyCompares_0_268;
  reg [3-1:0] put_KeyCollapse_0_269;
  reg [8-1:0] put_Data_0_270;
  reg [8-1:0] put_Key_1_271;
  reg [1-1:0] put_KeyCompares_1_272;
  reg [3-1:0] put_KeyCollapse_1_273;
  reg [8-1:0] put_Data_1_274;
  reg [8-1:0] put_Key_2_275;
  reg [1-1:0] put_KeyCompares_2_276;
  reg [3-1:0] put_KeyCollapse_2_277;
  reg [8-1:0] put_Data_2_278;
  reg [8-1:0] put_Key_3_279;
  reg [1-1:0] put_KeyCompares_3_280;
  reg [3-1:0] put_KeyCollapse_3_281;
  reg [8-1:0] put_Data_3_282;
  reg [1-1:0] put_Found_283;
  reg [8-1:0] put_Key_284;
  reg [8-1:0] put_FoundKey_285;
  reg [8-1:0] put_Data_286;
  reg [6-1:0] put_BtreeIndex_287;
  reg [3-1:0] put_StuckIndex_288;
  reg [1-1:0] put_MergeSuccess_289;
  reg [6-1:0] put_indexLeft_290;
  reg [6-1:0] put_indexRight_291;
  reg [8-1:0] put_midKey_292;
  reg [6-1:0] put_root_293;
  reg [6-1:0] put_next_294;
  reg [1-1:0] put_isLeaf_295;
  reg [1-1:0] put_isFree_296;
  reg [6-1:0] put_root_297;
  reg [6-1:0] put_next_298;
  reg [1-1:0] put_isLeaf_299;
  reg [1-1:0] put_isFree_300;
  reg [6-1:0] put_index_301;
  reg [3-1:0] put_size_302;
  reg [1-1:0] put_isLeaf_303;
  reg [6-1:0] put_nextFree_304;
  reg [8-1:0] put_Key_0_305;
  reg [1-1:0] put_KeyCompares_0_306;
  reg [3-1:0] put_KeyCollapse_0_307;
  reg [8-1:0] put_Data_0_308;
  reg [8-1:0] put_Key_1_309;
  reg [1-1:0] put_KeyCompares_1_310;
  reg [3-1:0] put_KeyCollapse_1_311;
  reg [8-1:0] put_Data_1_312;
  reg [8-1:0] put_Key_2_313;
  reg [1-1:0] put_KeyCompares_2_314;
  reg [3-1:0] put_KeyCollapse_2_315;
  reg [8-1:0] put_Data_2_316;
  reg [8-1:0] put_Key_3_317;
  reg [1-1:0] put_KeyCompares_3_318;
  reg [3-1:0] put_KeyCollapse_3_319;
  reg [8-1:0] put_Data_3_320;
  reg [1-1:0] put_Found_321;
  reg [8-1:0] put_Key_322;
  reg [8-1:0] put_FoundKey_323;
  reg [8-1:0] put_Data_324;
  reg [6-1:0] put_BtreeIndex_325;
  reg [3-1:0] put_StuckIndex_326;
  reg [1-1:0] put_MergeSuccess_327;
  reg [6-1:0] put_index_328;
  reg [3-1:0] put_size_329;
  reg [1-1:0] put_isLeaf_330;
  reg [6-1:0] put_nextFree_331;
  reg [8-1:0] put_Key_0_332;
  reg [1-1:0] put_KeyCompares_0_333;
  reg [3-1:0] put_KeyCollapse_0_334;
  reg [8-1:0] put_Data_0_335;
  reg [8-1:0] put_Key_1_336;
  reg [1-1:0] put_KeyCompares_1_337;
  reg [3-1:0] put_KeyCollapse_1_338;
  reg [8-1:0] put_Data_1_339;
  reg [8-1:0] put_Key_2_340;
  reg [1-1:0] put_KeyCompares_2_341;
  reg [3-1:0] put_KeyCollapse_2_342;
  reg [8-1:0] put_Data_2_343;
  reg [8-1:0] put_Key_3_344;
  reg [1-1:0] put_KeyCompares_3_345;
  reg [3-1:0] put_KeyCollapse_3_346;
  reg [8-1:0] put_Data_3_347;
  reg [1-1:0] put_Found_348;
  reg [8-1:0] put_Key_349;
  reg [8-1:0] put_FoundKey_350;
  reg [8-1:0] put_Data_351;
  reg [6-1:0] put_BtreeIndex_352;
  reg [3-1:0] put_StuckIndex_353;
  reg [1-1:0] put_MergeSuccess_354;
  reg [6-1:0] put_index_355;
  reg [3-1:0] put_size_356;
  reg [1-1:0] put_isLeaf_357;
  reg [6-1:0] put_nextFree_358;
  reg [8-1:0] put_Key_0_359;
  reg [1-1:0] put_KeyCompares_0_360;
  reg [3-1:0] put_KeyCollapse_0_361;
  reg [8-1:0] put_Data_0_362;
  reg [8-1:0] put_Key_1_363;
  reg [1-1:0] put_KeyCompares_1_364;
  reg [3-1:0] put_KeyCollapse_1_365;
  reg [8-1:0] put_Data_1_366;
  reg [8-1:0] put_Key_2_367;
  reg [1-1:0] put_KeyCompares_2_368;
  reg [3-1:0] put_KeyCollapse_2_369;
  reg [8-1:0] put_Data_2_370;
  reg [8-1:0] put_Key_3_371;
  reg [1-1:0] put_KeyCompares_3_372;
  reg [3-1:0] put_KeyCollapse_3_373;
  reg [8-1:0] put_Data_3_374;
  reg [1-1:0] put_Found_375;
  reg [8-1:0] put_Key_376;
  reg [8-1:0] put_FoundKey_377;
  reg [8-1:0] put_Data_378;
  reg [6-1:0] put_BtreeIndex_379;
  reg [3-1:0] put_StuckIndex_380;
  reg [1-1:0] put_MergeSuccess_381;
  reg [6-1:0] put_index_382;
  reg [3-1:0] put_size_383;
  reg [1-1:0] put_isLeaf_384;
  reg [6-1:0] put_nextFree_385;
  reg [8-1:0] put_Key_0_386;
  reg [1-1:0] put_KeyCompares_0_387;
  reg [3-1:0] put_KeyCollapse_0_388;
  reg [8-1:0] put_Data_0_389;
  reg [8-1:0] put_Key_1_390;
  reg [1-1:0] put_KeyCompares_1_391;
  reg [3-1:0] put_KeyCollapse_1_392;
  reg [8-1:0] put_Data_1_393;
  reg [8-1:0] put_Key_2_394;
  reg [1-1:0] put_KeyCompares_2_395;
  reg [3-1:0] put_KeyCollapse_2_396;
  reg [8-1:0] put_Data_2_397;
  reg [8-1:0] put_Key_3_398;
  reg [1-1:0] put_KeyCompares_3_399;
  reg [3-1:0] put_KeyCollapse_3_400;
  reg [8-1:0] put_Data_3_401;
  reg [1-1:0] put_Found_402;
  reg [8-1:0] put_Key_403;
  reg [8-1:0] put_FoundKey_404;
  reg [8-1:0] put_Data_405;
  reg [6-1:0] put_BtreeIndex_406;
  reg [3-1:0] put_StuckIndex_407;
  reg [1-1:0] put_MergeSuccess_408;
  reg [8-1:0] put_childKey_409;
  reg [6-1:0] put_childData_410;
  reg [6-1:0] put_indexLeft_411;
  reg [6-1:0] put_indexRight_412;
  reg [8-1:0] put_midKey_413;
  reg [6-1:0] put_root_414;
  reg [6-1:0] put_next_415;
  reg [1-1:0] put_isLeaf_416;
  reg [1-1:0] put_isFree_417;
  reg [6-1:0] put_index_418;
  reg [3-1:0] put_size_419;
  reg [1-1:0] put_isLeaf_420;
  reg [6-1:0] put_nextFree_421;
  reg [8-1:0] put_Key_0_422;
  reg [1-1:0] put_KeyCompares_0_423;
  reg [3-1:0] put_KeyCollapse_0_424;
  reg [8-1:0] put_Data_0_425;
  reg [8-1:0] put_Key_1_426;
  reg [1-1:0] put_KeyCompares_1_427;
  reg [3-1:0] put_KeyCollapse_1_428;
  reg [8-1:0] put_Data_1_429;
  reg [8-1:0] put_Key_2_430;
  reg [1-1:0] put_KeyCompares_2_431;
  reg [3-1:0] put_KeyCollapse_2_432;
  reg [8-1:0] put_Data_2_433;
  reg [8-1:0] put_Key_3_434;
  reg [1-1:0] put_KeyCompares_3_435;
  reg [3-1:0] put_KeyCollapse_3_436;
  reg [8-1:0] put_Data_3_437;
  reg [1-1:0] put_Found_438;
  reg [8-1:0] put_Key_439;
  reg [8-1:0] put_FoundKey_440;
  reg [8-1:0] put_Data_441;
  reg [6-1:0] put_BtreeIndex_442;
  reg [3-1:0] put_StuckIndex_443;
  reg [1-1:0] put_MergeSuccess_444;
  reg [6-1:0] put_index_445;
  reg [3-1:0] put_size_446;
  reg [1-1:0] put_isLeaf_447;
  reg [6-1:0] put_nextFree_448;
  reg [8-1:0] put_Key_0_449;
  reg [1-1:0] put_KeyCompares_0_450;
  reg [3-1:0] put_KeyCollapse_0_451;
  reg [8-1:0] put_Data_0_452;
  reg [8-1:0] put_Key_1_453;
  reg [1-1:0] put_KeyCompares_1_454;
  reg [3-1:0] put_KeyCollapse_1_455;
  reg [8-1:0] put_Data_1_456;
  reg [8-1:0] put_Key_2_457;
  reg [1-1:0] put_KeyCompares_2_458;
  reg [3-1:0] put_KeyCollapse_2_459;
  reg [8-1:0] put_Data_2_460;
  reg [8-1:0] put_Key_3_461;
  reg [1-1:0] put_KeyCompares_3_462;
  reg [3-1:0] put_KeyCollapse_3_463;
  reg [8-1:0] put_Data_3_464;
  reg [1-1:0] put_Found_465;
  reg [8-1:0] put_Key_466;
  reg [8-1:0] put_FoundKey_467;
  reg [8-1:0] put_Data_468;
  reg [6-1:0] put_BtreeIndex_469;
  reg [3-1:0] put_StuckIndex_470;
  reg [1-1:0] put_MergeSuccess_471;
  reg [6-1:0] put_index_472;
  reg [3-1:0] put_size_473;
  reg [1-1:0] put_isLeaf_474;
  reg [6-1:0] put_nextFree_475;
  reg [8-1:0] put_Key_0_476;
  reg [1-1:0] put_KeyCompares_0_477;
  reg [3-1:0] put_KeyCollapse_0_478;
  reg [8-1:0] put_Data_0_479;
  reg [8-1:0] put_Key_1_480;
  reg [1-1:0] put_KeyCompares_1_481;
  reg [3-1:0] put_KeyCollapse_1_482;
  reg [8-1:0] put_Data_1_483;
  reg [8-1:0] put_Key_2_484;
  reg [1-1:0] put_KeyCompares_2_485;
  reg [3-1:0] put_KeyCollapse_2_486;
  reg [8-1:0] put_Data_2_487;
  reg [8-1:0] put_Key_3_488;
  reg [1-1:0] put_KeyCompares_3_489;
  reg [3-1:0] put_KeyCollapse_3_490;
  reg [8-1:0] put_Data_3_491;
  reg [1-1:0] put_Found_492;
  reg [8-1:0] put_Key_493;
  reg [8-1:0] put_FoundKey_494;
  reg [8-1:0] put_Data_495;
  reg [6-1:0] put_BtreeIndex_496;
  reg [3-1:0] put_StuckIndex_497;
  reg [1-1:0] put_MergeSuccess_498;
  reg [6-1:0] put_childIndex_499;
  reg [6-1:0] put_leftIndex_500;
  reg [8-1:0] put_midKey_501;
  reg [6-1:0] put_root_502;
  reg [6-1:0] put_next_503;
  reg [1-1:0] put_isLeaf_504;
  reg [1-1:0] put_isFree_505;
  reg [3-1:0] put_i_506;
  reg [1-1:0] put_notFull_507;
  reg [6-1:0] put_index_508;
  reg [3-1:0] put_size_509;
  reg [1-1:0] put_isLeaf_510;
  reg [6-1:0] put_nextFree_511;
  reg [8-1:0] put_Key_0_512;
  reg [1-1:0] put_KeyCompares_0_513;
  reg [3-1:0] put_KeyCollapse_0_514;
  reg [8-1:0] put_Data_0_515;
  reg [8-1:0] put_Key_1_516;
  reg [1-1:0] put_KeyCompares_1_517;
  reg [3-1:0] put_KeyCollapse_1_518;
  reg [8-1:0] put_Data_1_519;
  reg [8-1:0] put_Key_2_520;
  reg [1-1:0] put_KeyCompares_2_521;
  reg [3-1:0] put_KeyCollapse_2_522;
  reg [8-1:0] put_Data_2_523;
  reg [8-1:0] put_Key_3_524;
  reg [1-1:0] put_KeyCompares_3_525;
  reg [3-1:0] put_KeyCollapse_3_526;
  reg [8-1:0] put_Data_3_527;
  reg [1-1:0] put_Found_528;
  reg [8-1:0] put_Key_529;
  reg [8-1:0] put_FoundKey_530;
  reg [8-1:0] put_Data_531;
  reg [6-1:0] put_BtreeIndex_532;
  reg [3-1:0] put_StuckIndex_533;
  reg [1-1:0] put_MergeSuccess_534;
  reg [6-1:0] put_index_535;
  reg [3-1:0] put_size_536;
  reg [1-1:0] put_isLeaf_537;
  reg [6-1:0] put_nextFree_538;
  reg [8-1:0] put_Key_0_539;
  reg [1-1:0] put_KeyCompares_0_540;
  reg [3-1:0] put_KeyCollapse_0_541;
  reg [8-1:0] put_Data_0_542;
  reg [8-1:0] put_Key_1_543;
  reg [1-1:0] put_KeyCompares_1_544;
  reg [3-1:0] put_KeyCollapse_1_545;
  reg [8-1:0] put_Data_1_546;
  reg [8-1:0] put_Key_2_547;
  reg [1-1:0] put_KeyCompares_2_548;
  reg [3-1:0] put_KeyCollapse_2_549;
  reg [8-1:0] put_Data_2_550;
  reg [8-1:0] put_Key_3_551;
  reg [1-1:0] put_KeyCompares_3_552;
  reg [3-1:0] put_KeyCollapse_3_553;
  reg [8-1:0] put_Data_3_554;
  reg [1-1:0] put_Found_555;
  reg [8-1:0] put_Key_556;
  reg [8-1:0] put_FoundKey_557;
  reg [8-1:0] put_Data_558;
  reg [6-1:0] put_BtreeIndex_559;
  reg [3-1:0] put_StuckIndex_560;
  reg [1-1:0] put_MergeSuccess_561;
  reg [6-1:0] put_index_562;
  reg [3-1:0] put_size_563;
  reg [1-1:0] put_isLeaf_564;
  reg [6-1:0] put_nextFree_565;
  reg [8-1:0] put_Key_0_566;
  reg [1-1:0] put_KeyCompares_0_567;
  reg [3-1:0] put_KeyCollapse_0_568;
  reg [8-1:0] put_Data_0_569;
  reg [8-1:0] put_Key_1_570;
  reg [1-1:0] put_KeyCompares_1_571;
  reg [3-1:0] put_KeyCollapse_1_572;
  reg [8-1:0] put_Data_1_573;
  reg [8-1:0] put_Key_2_574;
  reg [1-1:0] put_KeyCompares_2_575;
  reg [3-1:0] put_KeyCollapse_2_576;
  reg [8-1:0] put_Data_2_577;
  reg [8-1:0] put_Key_3_578;
  reg [1-1:0] put_KeyCompares_3_579;
  reg [3-1:0] put_KeyCollapse_3_580;
  reg [8-1:0] put_Data_3_581;
  reg [1-1:0] put_Found_582;
  reg [8-1:0] put_Key_583;
  reg [8-1:0] put_FoundKey_584;
  reg [8-1:0] put_Data_585;
  reg [6-1:0] put_BtreeIndex_586;
  reg [3-1:0] put_StuckIndex_587;
  reg [1-1:0] put_MergeSuccess_588;
  reg [6-1:0] put_index_589;
  reg [3-1:0] put_size_590;
  reg [1-1:0] put_isLeaf_591;
  reg [6-1:0] put_nextFree_592;
  reg [8-1:0] put_Key_0_593;
  reg [1-1:0] put_KeyCompares_0_594;
  reg [3-1:0] put_KeyCollapse_0_595;
  reg [8-1:0] put_Data_0_596;
  reg [8-1:0] put_Key_1_597;
  reg [1-1:0] put_KeyCompares_1_598;
  reg [3-1:0] put_KeyCollapse_1_599;
  reg [8-1:0] put_Data_1_600;
  reg [8-1:0] put_Key_2_601;
  reg [1-1:0] put_KeyCompares_2_602;
  reg [3-1:0] put_KeyCollapse_2_603;
  reg [8-1:0] put_Data_2_604;
  reg [8-1:0] put_Key_3_605;
  reg [1-1:0] put_KeyCompares_3_606;
  reg [3-1:0] put_KeyCollapse_3_607;
  reg [8-1:0] put_Data_3_608;
  reg [1-1:0] put_Found_609;
  reg [8-1:0] put_Key_610;
  reg [8-1:0] put_FoundKey_611;
  reg [8-1:0] put_Data_612;
  reg [6-1:0] put_BtreeIndex_613;
  reg [3-1:0] put_StuckIndex_614;
  reg [1-1:0] put_MergeSuccess_615;
  reg [8-1:0] put_childKey_616;
  reg [6-1:0] put_childData_617;
  reg [6-1:0] put_indexLeft_618;
  reg [6-1:0] put_indexRight_619;
  reg [8-1:0] put_midKey_620;
  reg [6-1:0] put_root_621;
  reg [6-1:0] put_next_622;
  reg [1-1:0] put_isLeaf_623;
  reg [1-1:0] put_isFree_624;
  reg [6-1:0] put_index_625;
  reg [3-1:0] put_size_626;
  reg [1-1:0] put_isLeaf_627;
  reg [6-1:0] put_nextFree_628;
  reg [8-1:0] put_Key_0_629;
  reg [1-1:0] put_KeyCompares_0_630;
  reg [3-1:0] put_KeyCollapse_0_631;
  reg [8-1:0] put_Data_0_632;
  reg [8-1:0] put_Key_1_633;
  reg [1-1:0] put_KeyCompares_1_634;
  reg [3-1:0] put_KeyCollapse_1_635;
  reg [8-1:0] put_Data_1_636;
  reg [8-1:0] put_Key_2_637;
  reg [1-1:0] put_KeyCompares_2_638;
  reg [3-1:0] put_KeyCollapse_2_639;
  reg [8-1:0] put_Data_2_640;
  reg [8-1:0] put_Key_3_641;
  reg [1-1:0] put_KeyCompares_3_642;
  reg [3-1:0] put_KeyCollapse_3_643;
  reg [8-1:0] put_Data_3_644;
  reg [1-1:0] put_Found_645;
  reg [8-1:0] put_Key_646;
  reg [8-1:0] put_FoundKey_647;
  reg [8-1:0] put_Data_648;
  reg [6-1:0] put_BtreeIndex_649;
  reg [3-1:0] put_StuckIndex_650;
  reg [1-1:0] put_MergeSuccess_651;
  reg [6-1:0] put_index_652;
  reg [3-1:0] put_size_653;
  reg [1-1:0] put_isLeaf_654;
  reg [6-1:0] put_nextFree_655;
  reg [8-1:0] put_Key_0_656;
  reg [1-1:0] put_KeyCompares_0_657;
  reg [3-1:0] put_KeyCollapse_0_658;
  reg [8-1:0] put_Data_0_659;
  reg [8-1:0] put_Key_1_660;
  reg [1-1:0] put_KeyCompares_1_661;
  reg [3-1:0] put_KeyCollapse_1_662;
  reg [8-1:0] put_Data_1_663;
  reg [8-1:0] put_Key_2_664;
  reg [1-1:0] put_KeyCompares_2_665;
  reg [3-1:0] put_KeyCollapse_2_666;
  reg [8-1:0] put_Data_2_667;
  reg [8-1:0] put_Key_3_668;
  reg [1-1:0] put_KeyCompares_3_669;
  reg [3-1:0] put_KeyCollapse_3_670;
  reg [8-1:0] put_Data_3_671;
  reg [1-1:0] put_Found_672;
  reg [8-1:0] put_Key_673;
  reg [8-1:0] put_FoundKey_674;
  reg [8-1:0] put_Data_675;
  reg [6-1:0] put_BtreeIndex_676;
  reg [3-1:0] put_StuckIndex_677;
  reg [1-1:0] put_MergeSuccess_678;
  reg [6-1:0] put_index_679;
  reg [3-1:0] put_size_680;
  reg [1-1:0] put_isLeaf_681;
  reg [6-1:0] put_nextFree_682;
  reg [8-1:0] put_Key_0_683;
  reg [1-1:0] put_KeyCompares_0_684;
  reg [3-1:0] put_KeyCollapse_0_685;
  reg [8-1:0] put_Data_0_686;
  reg [8-1:0] put_Key_1_687;
  reg [1-1:0] put_KeyCompares_1_688;
  reg [3-1:0] put_KeyCollapse_1_689;
  reg [8-1:0] put_Data_1_690;
  reg [8-1:0] put_Key_2_691;
  reg [1-1:0] put_KeyCompares_2_692;
  reg [3-1:0] put_KeyCollapse_2_693;
  reg [8-1:0] put_Data_2_694;
  reg [8-1:0] put_Key_3_695;
  reg [1-1:0] put_KeyCompares_3_696;
  reg [3-1:0] put_KeyCollapse_3_697;
  reg [8-1:0] put_Data_3_698;
  reg [1-1:0] put_Found_699;
  reg [8-1:0] put_Key_700;
  reg [8-1:0] put_FoundKey_701;
  reg [8-1:0] put_Data_702;
  reg [6-1:0] put_BtreeIndex_703;
  reg [3-1:0] put_StuckIndex_704;
  reg [1-1:0] put_MergeSuccess_705;
  reg [6-1:0] put_index_706;
  reg [3-1:0] put_size_707;
  reg [1-1:0] put_isLeaf_708;
  reg [6-1:0] put_nextFree_709;
  reg [8-1:0] put_Key_0_710;
  reg [1-1:0] put_KeyCompares_0_711;
  reg [3-1:0] put_KeyCollapse_0_712;
  reg [8-1:0] put_Data_0_713;
  reg [8-1:0] put_Key_1_714;
  reg [1-1:0] put_KeyCompares_1_715;
  reg [3-1:0] put_KeyCollapse_1_716;
  reg [8-1:0] put_Data_1_717;
  reg [8-1:0] put_Key_2_718;
  reg [1-1:0] put_KeyCompares_2_719;
  reg [3-1:0] put_KeyCollapse_2_720;
  reg [8-1:0] put_Data_2_721;
  reg [8-1:0] put_Key_3_722;
  reg [1-1:0] put_KeyCompares_3_723;
  reg [3-1:0] put_KeyCollapse_3_724;
  reg [8-1:0] put_Data_3_725;
  reg [1-1:0] put_Found_726;
  reg [8-1:0] put_Key_727;
  reg [8-1:0] put_FoundKey_728;
  reg [8-1:0] put_Data_729;
  reg [6-1:0] put_BtreeIndex_730;
  reg [3-1:0] put_StuckIndex_731;
  reg [1-1:0] put_MergeSuccess_732;
  reg [8-1:0] put_childKey_733;
  reg [6-1:0] put_childData_734;
  reg [6-1:0] put_indexLeft_735;
  reg [6-1:0] put_indexRight_736;
  reg [8-1:0] put_midKey_737;
  reg [6-1:0] put_root_738;
  reg [6-1:0] put_next_739;
  reg [1-1:0] put_isLeaf_740;
  reg [1-1:0] put_isFree_741;
  integer put_pc;
  integer put_stop;
  integer put_returnCode;
  always @ (posedge clock) begin
    if (step < 0) begin
      put_pc <= 0;
      put_stop <= 0;
      put_returnCode <= 0;
      put_k_0 <= 0;
      put_d_1 <= 0;
      put_i_2 <= 0;
      put_l_3 <= 0;
      put_index_4 <= 0;
      put_size_5 <= 0;
      put_isLeaf_6 <= 0;
      put_nextFree_7 <= 0;
      put_Key_0_8 <= 0;
      put_KeyCompares_0_9 <= 0;
      put_KeyCollapse_0_10 <= 0;
      put_Data_0_11 <= 0;
      put_Key_1_12 <= 0;
      put_KeyCompares_1_13 <= 0;
      put_KeyCollapse_1_14 <= 0;
      put_Data_1_15 <= 0;
      put_Key_2_16 <= 0;
      put_KeyCompares_2_17 <= 0;
      put_KeyCollapse_2_18 <= 0;
      put_Data_2_19 <= 0;
      put_Key_3_20 <= 0;
      put_KeyCompares_3_21 <= 0;
      put_KeyCollapse_3_22 <= 0;
      put_Data_3_23 <= 0;
      put_stuckKeys_1_index_24 <= 0;
      put_stuckKeys_2_index_25 <= 0;
      put_stuckKeys_2_value_26 <= 0;
      put_stuckKeys_2_value_27 <= 0;
      put_stuckKeys_2_value_28 <= 0;
      put_stuckKeys_2_value_29 <= 0;
      put_stuckData_3_index_30 <= 0;
      put_stuckData_4_index_31 <= 0;
      put_stuckData_4_value_32 <= 0;
      put_stuckData_4_value_33 <= 0;
      put_stuckData_4_value_34 <= 0;
      put_stuckData_4_value_35 <= 0;
      put_stuckSize_5_index_36 <= 0;
      put_stuckSize_6_index_37 <= 0;
      put_stuckSize_6_value_38 <= 0;
      put_stuckIsLeaf_7_index_39 <= 0;
      put_stuckIsLeaf_8_index_40 <= 0;
      put_stuckIsLeaf_8_value_41 <= 0;
      put_Found_42 <= 0;
      put_Key_43 <= 0;
      put_FoundKey_44 <= 0;
      put_Data_45 <= 0;
      put_BtreeIndex_46 <= 0;
      put_StuckIndex_47 <= 0;
      put_MergeSuccess_48 <= 0;
      put_index_49 <= 0;
      put_size_50 <= 0;
      put_isLeaf_51 <= 0;
      put_nextFree_52 <= 0;
      put_Key_0_53 <= 0;
      put_KeyCompares_0_54 <= 0;
      put_KeyCollapse_0_55 <= 0;
      put_Data_0_56 <= 0;
      put_Key_1_57 <= 0;
      put_KeyCompares_1_58 <= 0;
      put_KeyCollapse_1_59 <= 0;
      put_Data_1_60 <= 0;
      put_Key_2_61 <= 0;
      put_KeyCompares_2_62 <= 0;
      put_KeyCollapse_2_63 <= 0;
      put_Data_2_64 <= 0;
      put_Key_3_65 <= 0;
      put_KeyCompares_3_66 <= 0;
      put_KeyCollapse_3_67 <= 0;
      put_Data_3_68 <= 0;
      put_Found_69 <= 0;
      put_Key_70 <= 0;
      put_FoundKey_71 <= 0;
      put_Data_72 <= 0;
      put_BtreeIndex_73 <= 0;
      put_StuckIndex_74 <= 0;
      put_MergeSuccess_75 <= 0;
      put_index_76 <= 0;
      put_size_77 <= 0;
      put_isLeaf_78 <= 0;
      put_nextFree_79 <= 0;
      put_Key_0_80 <= 0;
      put_KeyCompares_0_81 <= 0;
      put_KeyCollapse_0_82 <= 0;
      put_Data_0_83 <= 0;
      put_Key_1_84 <= 0;
      put_KeyCompares_1_85 <= 0;
      put_KeyCollapse_1_86 <= 0;
      put_Data_1_87 <= 0;
      put_Key_2_88 <= 0;
      put_KeyCompares_2_89 <= 0;
      put_KeyCollapse_2_90 <= 0;
      put_Data_2_91 <= 0;
      put_Key_3_92 <= 0;
      put_KeyCompares_3_93 <= 0;
      put_KeyCollapse_3_94 <= 0;
      put_Data_3_95 <= 0;
      put_Found_96 <= 0;
      put_Key_97 <= 0;
      put_FoundKey_98 <= 0;
      put_Data_99 <= 0;
      put_BtreeIndex_100 <= 0;
      put_StuckIndex_101 <= 0;
      put_MergeSuccess_102 <= 0;
      put_child_103 <= 0;
      put_parent_104 <= 0;
      put_childInparent_105 <= 0;
      put_found_106 <= 0;
      put_full_107 <= 0;
      put_i_108 <= 0;
      put_notFull_109 <= 0;
      put_index_110 <= 0;
      put_size_111 <= 0;
      put_isLeaf_112 <= 0;
      put_nextFree_113 <= 0;
      put_Key_0_114 <= 0;
      put_KeyCompares_0_115 <= 0;
      put_KeyCollapse_0_116 <= 0;
      put_Data_0_117 <= 0;
      put_Key_1_118 <= 0;
      put_KeyCompares_1_119 <= 0;
      put_KeyCollapse_1_120 <= 0;
      put_Data_1_121 <= 0;
      put_Key_2_122 <= 0;
      put_KeyCompares_2_123 <= 0;
      put_KeyCollapse_2_124 <= 0;
      put_Data_2_125 <= 0;
      put_Key_3_126 <= 0;
      put_KeyCompares_3_127 <= 0;
      put_KeyCollapse_3_128 <= 0;
      put_Data_3_129 <= 0;
      put_Found_130 <= 0;
      put_Key_131 <= 0;
      put_FoundKey_132 <= 0;
      put_Data_133 <= 0;
      put_BtreeIndex_134 <= 0;
      put_StuckIndex_135 <= 0;
      put_MergeSuccess_136 <= 0;
      put_index_137 <= 0;
      put_size_138 <= 0;
      put_isLeaf_139 <= 0;
      put_nextFree_140 <= 0;
      put_Key_0_141 <= 0;
      put_KeyCompares_0_142 <= 0;
      put_KeyCollapse_0_143 <= 0;
      put_Data_0_144 <= 0;
      put_Key_1_145 <= 0;
      put_KeyCompares_1_146 <= 0;
      put_KeyCollapse_1_147 <= 0;
      put_Data_1_148 <= 0;
      put_Key_2_149 <= 0;
      put_KeyCompares_2_150 <= 0;
      put_KeyCollapse_2_151 <= 0;
      put_Data_2_152 <= 0;
      put_Key_3_153 <= 0;
      put_KeyCompares_3_154 <= 0;
      put_KeyCollapse_3_155 <= 0;
      put_Data_3_156 <= 0;
      put_Found_157 <= 0;
      put_Key_158 <= 0;
      put_FoundKey_159 <= 0;
      put_Data_160 <= 0;
      put_BtreeIndex_161 <= 0;
      put_StuckIndex_162 <= 0;
      put_MergeSuccess_163 <= 0;
      put_index_164 <= 0;
      put_size_165 <= 0;
      put_isLeaf_166 <= 0;
      put_nextFree_167 <= 0;
      put_Key_0_168 <= 0;
      put_KeyCompares_0_169 <= 0;
      put_KeyCollapse_0_170 <= 0;
      put_Data_0_171 <= 0;
      put_Key_1_172 <= 0;
      put_KeyCompares_1_173 <= 0;
      put_KeyCollapse_1_174 <= 0;
      put_Data_1_175 <= 0;
      put_Key_2_176 <= 0;
      put_KeyCompares_2_177 <= 0;
      put_KeyCollapse_2_178 <= 0;
      put_Data_2_179 <= 0;
      put_Key_3_180 <= 0;
      put_KeyCompares_3_181 <= 0;
      put_KeyCollapse_3_182 <= 0;
      put_Data_3_183 <= 0;
      put_Found_184 <= 0;
      put_Key_185 <= 0;
      put_FoundKey_186 <= 0;
      put_Data_187 <= 0;
      put_BtreeIndex_188 <= 0;
      put_StuckIndex_189 <= 0;
      put_MergeSuccess_190 <= 0;
      put_indexLeft_191 <= 0;
      put_indexRight_192 <= 0;
      put_midKey_193 <= 0;
      put_freeNext_9_index_194 <= 0;
      put_freeNext_10_index_195 <= 0;
      put_freeNext_10_value_196 <= 0;
      put_stuckIsFree_11_index_197 <= 0;
      put_stuckIsFree_11_value_198 <= 0;
      put_root_199 <= 0;
      put_next_200 <= 0;
      put_isLeaf_201 <= 0;
      put_isFree_202 <= 0;
      put_root_203 <= 0;
      put_next_204 <= 0;
      put_isLeaf_205 <= 0;
      put_isFree_206 <= 0;
      put_i_207 <= 0;
      put_notFull_208 <= 0;
      put_index_209 <= 0;
      put_size_210 <= 0;
      put_isLeaf_211 <= 0;
      put_nextFree_212 <= 0;
      put_Key_0_213 <= 0;
      put_KeyCompares_0_214 <= 0;
      put_KeyCollapse_0_215 <= 0;
      put_Data_0_216 <= 0;
      put_Key_1_217 <= 0;
      put_KeyCompares_1_218 <= 0;
      put_KeyCollapse_1_219 <= 0;
      put_Data_1_220 <= 0;
      put_Key_2_221 <= 0;
      put_KeyCompares_2_222 <= 0;
      put_KeyCollapse_2_223 <= 0;
      put_Data_2_224 <= 0;
      put_Key_3_225 <= 0;
      put_KeyCompares_3_226 <= 0;
      put_KeyCollapse_3_227 <= 0;
      put_Data_3_228 <= 0;
      put_Found_229 <= 0;
      put_Key_230 <= 0;
      put_FoundKey_231 <= 0;
      put_Data_232 <= 0;
      put_BtreeIndex_233 <= 0;
      put_StuckIndex_234 <= 0;
      put_MergeSuccess_235 <= 0;
      put_index_236 <= 0;
      put_size_237 <= 0;
      put_isLeaf_238 <= 0;
      put_nextFree_239 <= 0;
      put_Key_0_240 <= 0;
      put_KeyCompares_0_241 <= 0;
      put_KeyCollapse_0_242 <= 0;
      put_Data_0_243 <= 0;
      put_Key_1_244 <= 0;
      put_KeyCompares_1_245 <= 0;
      put_KeyCollapse_1_246 <= 0;
      put_Data_1_247 <= 0;
      put_Key_2_248 <= 0;
      put_KeyCompares_2_249 <= 0;
      put_KeyCollapse_2_250 <= 0;
      put_Data_2_251 <= 0;
      put_Key_3_252 <= 0;
      put_KeyCompares_3_253 <= 0;
      put_KeyCollapse_3_254 <= 0;
      put_Data_3_255 <= 0;
      put_Found_256 <= 0;
      put_Key_257 <= 0;
      put_FoundKey_258 <= 0;
      put_Data_259 <= 0;
      put_BtreeIndex_260 <= 0;
      put_StuckIndex_261 <= 0;
      put_MergeSuccess_262 <= 0;
      put_index_263 <= 0;
      put_size_264 <= 0;
      put_isLeaf_265 <= 0;
      put_nextFree_266 <= 0;
      put_Key_0_267 <= 0;
      put_KeyCompares_0_268 <= 0;
      put_KeyCollapse_0_269 <= 0;
      put_Data_0_270 <= 0;
      put_Key_1_271 <= 0;
      put_KeyCompares_1_272 <= 0;
      put_KeyCollapse_1_273 <= 0;
      put_Data_1_274 <= 0;
      put_Key_2_275 <= 0;
      put_KeyCompares_2_276 <= 0;
      put_KeyCollapse_2_277 <= 0;
      put_Data_2_278 <= 0;
      put_Key_3_279 <= 0;
      put_KeyCompares_3_280 <= 0;
      put_KeyCollapse_3_281 <= 0;
      put_Data_3_282 <= 0;
      put_Found_283 <= 0;
      put_Key_284 <= 0;
      put_FoundKey_285 <= 0;
      put_Data_286 <= 0;
      put_BtreeIndex_287 <= 0;
      put_StuckIndex_288 <= 0;
      put_MergeSuccess_289 <= 0;
      put_indexLeft_290 <= 0;
      put_indexRight_291 <= 0;
      put_midKey_292 <= 0;
      put_root_293 <= 0;
      put_next_294 <= 0;
      put_isLeaf_295 <= 0;
      put_isFree_296 <= 0;
      put_root_297 <= 0;
      put_next_298 <= 0;
      put_isLeaf_299 <= 0;
      put_isFree_300 <= 0;
      put_index_301 <= 0;
      put_size_302 <= 0;
      put_isLeaf_303 <= 0;
      put_nextFree_304 <= 0;
      put_Key_0_305 <= 0;
      put_KeyCompares_0_306 <= 0;
      put_KeyCollapse_0_307 <= 0;
      put_Data_0_308 <= 0;
      put_Key_1_309 <= 0;
      put_KeyCompares_1_310 <= 0;
      put_KeyCollapse_1_311 <= 0;
      put_Data_1_312 <= 0;
      put_Key_2_313 <= 0;
      put_KeyCompares_2_314 <= 0;
      put_KeyCollapse_2_315 <= 0;
      put_Data_2_316 <= 0;
      put_Key_3_317 <= 0;
      put_KeyCompares_3_318 <= 0;
      put_KeyCollapse_3_319 <= 0;
      put_Data_3_320 <= 0;
      put_Found_321 <= 0;
      put_Key_322 <= 0;
      put_FoundKey_323 <= 0;
      put_Data_324 <= 0;
      put_BtreeIndex_325 <= 0;
      put_StuckIndex_326 <= 0;
      put_MergeSuccess_327 <= 0;
      put_index_328 <= 0;
      put_size_329 <= 0;
      put_isLeaf_330 <= 0;
      put_nextFree_331 <= 0;
      put_Key_0_332 <= 0;
      put_KeyCompares_0_333 <= 0;
      put_KeyCollapse_0_334 <= 0;
      put_Data_0_335 <= 0;
      put_Key_1_336 <= 0;
      put_KeyCompares_1_337 <= 0;
      put_KeyCollapse_1_338 <= 0;
      put_Data_1_339 <= 0;
      put_Key_2_340 <= 0;
      put_KeyCompares_2_341 <= 0;
      put_KeyCollapse_2_342 <= 0;
      put_Data_2_343 <= 0;
      put_Key_3_344 <= 0;
      put_KeyCompares_3_345 <= 0;
      put_KeyCollapse_3_346 <= 0;
      put_Data_3_347 <= 0;
      put_Found_348 <= 0;
      put_Key_349 <= 0;
      put_FoundKey_350 <= 0;
      put_Data_351 <= 0;
      put_BtreeIndex_352 <= 0;
      put_StuckIndex_353 <= 0;
      put_MergeSuccess_354 <= 0;
      put_index_355 <= 0;
      put_size_356 <= 0;
      put_isLeaf_357 <= 0;
      put_nextFree_358 <= 0;
      put_Key_0_359 <= 0;
      put_KeyCompares_0_360 <= 0;
      put_KeyCollapse_0_361 <= 0;
      put_Data_0_362 <= 0;
      put_Key_1_363 <= 0;
      put_KeyCompares_1_364 <= 0;
      put_KeyCollapse_1_365 <= 0;
      put_Data_1_366 <= 0;
      put_Key_2_367 <= 0;
      put_KeyCompares_2_368 <= 0;
      put_KeyCollapse_2_369 <= 0;
      put_Data_2_370 <= 0;
      put_Key_3_371 <= 0;
      put_KeyCompares_3_372 <= 0;
      put_KeyCollapse_3_373 <= 0;
      put_Data_3_374 <= 0;
      put_Found_375 <= 0;
      put_Key_376 <= 0;
      put_FoundKey_377 <= 0;
      put_Data_378 <= 0;
      put_BtreeIndex_379 <= 0;
      put_StuckIndex_380 <= 0;
      put_MergeSuccess_381 <= 0;
      put_index_382 <= 0;
      put_size_383 <= 0;
      put_isLeaf_384 <= 0;
      put_nextFree_385 <= 0;
      put_Key_0_386 <= 0;
      put_KeyCompares_0_387 <= 0;
      put_KeyCollapse_0_388 <= 0;
      put_Data_0_389 <= 0;
      put_Key_1_390 <= 0;
      put_KeyCompares_1_391 <= 0;
      put_KeyCollapse_1_392 <= 0;
      put_Data_1_393 <= 0;
      put_Key_2_394 <= 0;
      put_KeyCompares_2_395 <= 0;
      put_KeyCollapse_2_396 <= 0;
      put_Data_2_397 <= 0;
      put_Key_3_398 <= 0;
      put_KeyCompares_3_399 <= 0;
      put_KeyCollapse_3_400 <= 0;
      put_Data_3_401 <= 0;
      put_Found_402 <= 0;
      put_Key_403 <= 0;
      put_FoundKey_404 <= 0;
      put_Data_405 <= 0;
      put_BtreeIndex_406 <= 0;
      put_StuckIndex_407 <= 0;
      put_MergeSuccess_408 <= 0;
      put_childKey_409 <= 0;
      put_childData_410 <= 0;
      put_indexLeft_411 <= 0;
      put_indexRight_412 <= 0;
      put_midKey_413 <= 0;
      put_root_414 <= 0;
      put_next_415 <= 0;
      put_isLeaf_416 <= 0;
      put_isFree_417 <= 0;
      put_index_418 <= 0;
      put_size_419 <= 0;
      put_isLeaf_420 <= 0;
      put_nextFree_421 <= 0;
      put_Key_0_422 <= 0;
      put_KeyCompares_0_423 <= 0;
      put_KeyCollapse_0_424 <= 0;
      put_Data_0_425 <= 0;
      put_Key_1_426 <= 0;
      put_KeyCompares_1_427 <= 0;
      put_KeyCollapse_1_428 <= 0;
      put_Data_1_429 <= 0;
      put_Key_2_430 <= 0;
      put_KeyCompares_2_431 <= 0;
      put_KeyCollapse_2_432 <= 0;
      put_Data_2_433 <= 0;
      put_Key_3_434 <= 0;
      put_KeyCompares_3_435 <= 0;
      put_KeyCollapse_3_436 <= 0;
      put_Data_3_437 <= 0;
      put_Found_438 <= 0;
      put_Key_439 <= 0;
      put_FoundKey_440 <= 0;
      put_Data_441 <= 0;
      put_BtreeIndex_442 <= 0;
      put_StuckIndex_443 <= 0;
      put_MergeSuccess_444 <= 0;
      put_index_445 <= 0;
      put_size_446 <= 0;
      put_isLeaf_447 <= 0;
      put_nextFree_448 <= 0;
      put_Key_0_449 <= 0;
      put_KeyCompares_0_450 <= 0;
      put_KeyCollapse_0_451 <= 0;
      put_Data_0_452 <= 0;
      put_Key_1_453 <= 0;
      put_KeyCompares_1_454 <= 0;
      put_KeyCollapse_1_455 <= 0;
      put_Data_1_456 <= 0;
      put_Key_2_457 <= 0;
      put_KeyCompares_2_458 <= 0;
      put_KeyCollapse_2_459 <= 0;
      put_Data_2_460 <= 0;
      put_Key_3_461 <= 0;
      put_KeyCompares_3_462 <= 0;
      put_KeyCollapse_3_463 <= 0;
      put_Data_3_464 <= 0;
      put_Found_465 <= 0;
      put_Key_466 <= 0;
      put_FoundKey_467 <= 0;
      put_Data_468 <= 0;
      put_BtreeIndex_469 <= 0;
      put_StuckIndex_470 <= 0;
      put_MergeSuccess_471 <= 0;
      put_index_472 <= 0;
      put_size_473 <= 0;
      put_isLeaf_474 <= 0;
      put_nextFree_475 <= 0;
      put_Key_0_476 <= 0;
      put_KeyCompares_0_477 <= 0;
      put_KeyCollapse_0_478 <= 0;
      put_Data_0_479 <= 0;
      put_Key_1_480 <= 0;
      put_KeyCompares_1_481 <= 0;
      put_KeyCollapse_1_482 <= 0;
      put_Data_1_483 <= 0;
      put_Key_2_484 <= 0;
      put_KeyCompares_2_485 <= 0;
      put_KeyCollapse_2_486 <= 0;
      put_Data_2_487 <= 0;
      put_Key_3_488 <= 0;
      put_KeyCompares_3_489 <= 0;
      put_KeyCollapse_3_490 <= 0;
      put_Data_3_491 <= 0;
      put_Found_492 <= 0;
      put_Key_493 <= 0;
      put_FoundKey_494 <= 0;
      put_Data_495 <= 0;
      put_BtreeIndex_496 <= 0;
      put_StuckIndex_497 <= 0;
      put_MergeSuccess_498 <= 0;
      put_childIndex_499 <= 0;
      put_leftIndex_500 <= 0;
      put_midKey_501 <= 0;
      put_root_502 <= 0;
      put_next_503 <= 0;
      put_isLeaf_504 <= 0;
      put_isFree_505 <= 0;
      put_i_506 <= 0;
      put_notFull_507 <= 0;
      put_index_508 <= 0;
      put_size_509 <= 0;
      put_isLeaf_510 <= 0;
      put_nextFree_511 <= 0;
      put_Key_0_512 <= 0;
      put_KeyCompares_0_513 <= 0;
      put_KeyCollapse_0_514 <= 0;
      put_Data_0_515 <= 0;
      put_Key_1_516 <= 0;
      put_KeyCompares_1_517 <= 0;
      put_KeyCollapse_1_518 <= 0;
      put_Data_1_519 <= 0;
      put_Key_2_520 <= 0;
      put_KeyCompares_2_521 <= 0;
      put_KeyCollapse_2_522 <= 0;
      put_Data_2_523 <= 0;
      put_Key_3_524 <= 0;
      put_KeyCompares_3_525 <= 0;
      put_KeyCollapse_3_526 <= 0;
      put_Data_3_527 <= 0;
      put_Found_528 <= 0;
      put_Key_529 <= 0;
      put_FoundKey_530 <= 0;
      put_Data_531 <= 0;
      put_BtreeIndex_532 <= 0;
      put_StuckIndex_533 <= 0;
      put_MergeSuccess_534 <= 0;
      put_index_535 <= 0;
      put_size_536 <= 0;
      put_isLeaf_537 <= 0;
      put_nextFree_538 <= 0;
      put_Key_0_539 <= 0;
      put_KeyCompares_0_540 <= 0;
      put_KeyCollapse_0_541 <= 0;
      put_Data_0_542 <= 0;
      put_Key_1_543 <= 0;
      put_KeyCompares_1_544 <= 0;
      put_KeyCollapse_1_545 <= 0;
      put_Data_1_546 <= 0;
      put_Key_2_547 <= 0;
      put_KeyCompares_2_548 <= 0;
      put_KeyCollapse_2_549 <= 0;
      put_Data_2_550 <= 0;
      put_Key_3_551 <= 0;
      put_KeyCompares_3_552 <= 0;
      put_KeyCollapse_3_553 <= 0;
      put_Data_3_554 <= 0;
      put_Found_555 <= 0;
      put_Key_556 <= 0;
      put_FoundKey_557 <= 0;
      put_Data_558 <= 0;
      put_BtreeIndex_559 <= 0;
      put_StuckIndex_560 <= 0;
      put_MergeSuccess_561 <= 0;
      put_index_562 <= 0;
      put_size_563 <= 0;
      put_isLeaf_564 <= 0;
      put_nextFree_565 <= 0;
      put_Key_0_566 <= 0;
      put_KeyCompares_0_567 <= 0;
      put_KeyCollapse_0_568 <= 0;
      put_Data_0_569 <= 0;
      put_Key_1_570 <= 0;
      put_KeyCompares_1_571 <= 0;
      put_KeyCollapse_1_572 <= 0;
      put_Data_1_573 <= 0;
      put_Key_2_574 <= 0;
      put_KeyCompares_2_575 <= 0;
      put_KeyCollapse_2_576 <= 0;
      put_Data_2_577 <= 0;
      put_Key_3_578 <= 0;
      put_KeyCompares_3_579 <= 0;
      put_KeyCollapse_3_580 <= 0;
      put_Data_3_581 <= 0;
      put_Found_582 <= 0;
      put_Key_583 <= 0;
      put_FoundKey_584 <= 0;
      put_Data_585 <= 0;
      put_BtreeIndex_586 <= 0;
      put_StuckIndex_587 <= 0;
      put_MergeSuccess_588 <= 0;
      put_index_589 <= 0;
      put_size_590 <= 0;
      put_isLeaf_591 <= 0;
      put_nextFree_592 <= 0;
      put_Key_0_593 <= 0;
      put_KeyCompares_0_594 <= 0;
      put_KeyCollapse_0_595 <= 0;
      put_Data_0_596 <= 0;
      put_Key_1_597 <= 0;
      put_KeyCompares_1_598 <= 0;
      put_KeyCollapse_1_599 <= 0;
      put_Data_1_600 <= 0;
      put_Key_2_601 <= 0;
      put_KeyCompares_2_602 <= 0;
      put_KeyCollapse_2_603 <= 0;
      put_Data_2_604 <= 0;
      put_Key_3_605 <= 0;
      put_KeyCompares_3_606 <= 0;
      put_KeyCollapse_3_607 <= 0;
      put_Data_3_608 <= 0;
      put_Found_609 <= 0;
      put_Key_610 <= 0;
      put_FoundKey_611 <= 0;
      put_Data_612 <= 0;
      put_BtreeIndex_613 <= 0;
      put_StuckIndex_614 <= 0;
      put_MergeSuccess_615 <= 0;
      put_childKey_616 <= 0;
      put_childData_617 <= 0;
      put_indexLeft_618 <= 0;
      put_indexRight_619 <= 0;
      put_midKey_620 <= 0;
      put_root_621 <= 0;
      put_next_622 <= 0;
      put_isLeaf_623 <= 0;
      put_isFree_624 <= 0;
      put_index_625 <= 0;
      put_size_626 <= 0;
      put_isLeaf_627 <= 0;
      put_nextFree_628 <= 0;
      put_Key_0_629 <= 0;
      put_KeyCompares_0_630 <= 0;
      put_KeyCollapse_0_631 <= 0;
      put_Data_0_632 <= 0;
      put_Key_1_633 <= 0;
      put_KeyCompares_1_634 <= 0;
      put_KeyCollapse_1_635 <= 0;
      put_Data_1_636 <= 0;
      put_Key_2_637 <= 0;
      put_KeyCompares_2_638 <= 0;
      put_KeyCollapse_2_639 <= 0;
      put_Data_2_640 <= 0;
      put_Key_3_641 <= 0;
      put_KeyCompares_3_642 <= 0;
      put_KeyCollapse_3_643 <= 0;
      put_Data_3_644 <= 0;
      put_Found_645 <= 0;
      put_Key_646 <= 0;
      put_FoundKey_647 <= 0;
      put_Data_648 <= 0;
      put_BtreeIndex_649 <= 0;
      put_StuckIndex_650 <= 0;
      put_MergeSuccess_651 <= 0;
      put_index_652 <= 0;
      put_size_653 <= 0;
      put_isLeaf_654 <= 0;
      put_nextFree_655 <= 0;
      put_Key_0_656 <= 0;
      put_KeyCompares_0_657 <= 0;
      put_KeyCollapse_0_658 <= 0;
      put_Data_0_659 <= 0;
      put_Key_1_660 <= 0;
      put_KeyCompares_1_661 <= 0;
      put_KeyCollapse_1_662 <= 0;
      put_Data_1_663 <= 0;
      put_Key_2_664 <= 0;
      put_KeyCompares_2_665 <= 0;
      put_KeyCollapse_2_666 <= 0;
      put_Data_2_667 <= 0;
      put_Key_3_668 <= 0;
      put_KeyCompares_3_669 <= 0;
      put_KeyCollapse_3_670 <= 0;
      put_Data_3_671 <= 0;
      put_Found_672 <= 0;
      put_Key_673 <= 0;
      put_FoundKey_674 <= 0;
      put_Data_675 <= 0;
      put_BtreeIndex_676 <= 0;
      put_StuckIndex_677 <= 0;
      put_MergeSuccess_678 <= 0;
      put_index_679 <= 0;
      put_size_680 <= 0;
      put_isLeaf_681 <= 0;
      put_nextFree_682 <= 0;
      put_Key_0_683 <= 0;
      put_KeyCompares_0_684 <= 0;
      put_KeyCollapse_0_685 <= 0;
      put_Data_0_686 <= 0;
      put_Key_1_687 <= 0;
      put_KeyCompares_1_688 <= 0;
      put_KeyCollapse_1_689 <= 0;
      put_Data_1_690 <= 0;
      put_Key_2_691 <= 0;
      put_KeyCompares_2_692 <= 0;
      put_KeyCollapse_2_693 <= 0;
      put_Data_2_694 <= 0;
      put_Key_3_695 <= 0;
      put_KeyCompares_3_696 <= 0;
      put_KeyCollapse_3_697 <= 0;
      put_Data_3_698 <= 0;
      put_Found_699 <= 0;
      put_Key_700 <= 0;
      put_FoundKey_701 <= 0;
      put_Data_702 <= 0;
      put_BtreeIndex_703 <= 0;
      put_StuckIndex_704 <= 0;
      put_MergeSuccess_705 <= 0;
      put_index_706 <= 0;
      put_size_707 <= 0;
      put_isLeaf_708 <= 0;
      put_nextFree_709 <= 0;
      put_Key_0_710 <= 0;
      put_KeyCompares_0_711 <= 0;
      put_KeyCollapse_0_712 <= 0;
      put_Data_0_713 <= 0;
      put_Key_1_714 <= 0;
      put_KeyCompares_1_715 <= 0;
      put_KeyCollapse_1_716 <= 0;
      put_Data_1_717 <= 0;
      put_Key_2_718 <= 0;
      put_KeyCompares_2_719 <= 0;
      put_KeyCollapse_2_720 <= 0;
      put_Data_2_721 <= 0;
      put_Key_3_722 <= 0;
      put_KeyCompares_3_723 <= 0;
      put_KeyCollapse_3_724 <= 0;
      put_Data_3_725 <= 0;
      put_Found_726 <= 0;
      put_Key_727 <= 0;
      put_FoundKey_728 <= 0;
      put_Data_729 <= 0;
      put_BtreeIndex_730 <= 0;
      put_StuckIndex_731 <= 0;
      put_MergeSuccess_732 <= 0;
      put_childKey_733 <= 0;
      put_childData_734 <= 0;
      put_indexLeft_735 <= 0;
      put_indexRight_736 <= 0;
      put_midKey_737 <= 0;
      put_root_738 <= 0;
      put_next_739 <= 0;
      put_isLeaf_740 <= 0;
      put_isFree_741 <= 0;
      stuckIsLeaf_7_requestedAt <= -1;
      stuckIsLeaf_8_requestedAt <= -1;
      stuckIsFree_11_requestedAt <= -1;
      freeNext_9_requestedAt <= -1;
      freeNext_10_requestedAt <= -1;
      stuckSize_5_requestedAt <= -1;
      stuckSize_6_requestedAt <= -1;
      stuckKeys_1_requestedAt <= -1;
      stuckKeys_2_requestedAt <= -1;
      stuckData_3_requestedAt <= -1;
      stuckData_4_requestedAt <= -1;
    end
    else if (processCurrent == 6) begin
      case(put_pc)
        0: begin
          put_k_0 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0676:<init>|  Chip.java:0675:RegisterSet|  Btree.java:5937:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        1: begin
          put_d_1 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0676:<init>|  Chip.java:0675:RegisterSet|  Btree.java:5938:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        2: begin
          put_k_0 <= put_k_0+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0806:<init>|  Chip.java:0805:Inc|  Btree.java:5941:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        3: begin
          put_d_1 <= put_k_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:5941:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        4: begin
          put_d_1 <= put_d_1+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0806:<init>|  Chip.java:0805:Inc|  Btree.java:5941:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        5: begin
          put_BtreeIndex_100 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        6: begin
          put_index_76 <= put_BtreeIndex_100;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        7: begin
          put_stuckSize_5_index_36 <= put_index_76;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_76;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_76;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_76;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        8: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        9: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        10: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        11: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        12: begin
          put_size_77 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_78 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_80 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_83 <= stuckData_stuckData_3_result_0;
          put_Key_1_84 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_87 <= stuckData_stuckData_3_result_1;
          put_Key_2_88 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_91 <= stuckData_stuckData_3_result_2;
          put_Key_3_92 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_95 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        13: begin
          if (put_isLeaf_78 == 0) begin
            put_pc <= 20;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1395:<init>|  Btree.java:1394:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        14: begin
          put_KeyCompares_0_81 <= put_k_0 == put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 == put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 == put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 == put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0802:<init>|  Btree.java:0801:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        15: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0823:<init>|  Btree.java:0822:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        16: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0823:<init>|  Btree.java:0822:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        17: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Key_97 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Key_97 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Key_97 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Key_97 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0845:<init>|  Btree.java:0844:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        18: begin
          put_pc <= 26;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2260:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        19: begin
          put_pc <= 26;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1411:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        20: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        21: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        22: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        23: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        24: begin
          put_BtreeIndex_100 <= put_Data_99;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2264:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        25: begin
          put_pc <= 6;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2265:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        26: begin
          if (put_Found_96 == 0) begin
            put_pc <= 29;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        27: begin
          if (put_StuckIndex_101 == put_size_77) begin
            put_size_77 <= put_size_77+1;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0626:<init>|  Btree.java:0625:SetElementAt|  Btree.java:2295:Then|  Chip.java:0610:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        28: begin
          put_pc <= 40;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        29: begin
          put_notFull_109 <= put_size_77< 4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        30: begin
          if (put_notFull_109 == 0) begin
            put_pc <= 39;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        31: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        32: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        33: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        34: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        35: begin
          put_size_77 <= put_size_77+1;
          if (3 > put_StuckIndex_101) begin
            put_Key_3_92 <= put_Key_2_88;
            put_Data_3_95 <= put_Data_2_91;
          end
          if (2 > put_StuckIndex_101) begin
            put_Key_2_88 <= put_Key_1_84;
            put_Data_2_91 <= put_Data_1_87;
          end
          if (1 > put_StuckIndex_101) begin
            put_Key_1_84 <= put_Key_0_80;
            put_Data_1_87 <= put_Data_0_83;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0701:<init>|  Btree.java:0700:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        36: begin
          put_Found_96 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2305:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        37: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0592:<init>|  Chip.java:0591:COntinue|  Btree.java:2306:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        38: begin
          put_pc <= 40;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        39: begin
          put_pc <= 44;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2309:Else|  Chip.java:0620:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        40: begin
          put_stuckSize_6_index_37 <= put_index_76;
          put_stuckSize_6_value_38 <= put_size_77;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_76;
          put_stuckKeys_2_value_26 <= put_Key_0_80;
          put_stuckKeys_2_value_27 <= put_Key_1_84;
          put_stuckKeys_2_value_28 <= put_Key_2_88;
          put_stuckKeys_2_value_29 <= put_Key_3_92;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_76;
          put_stuckData_4_value_32 <= put_Data_0_83;
          put_stuckData_4_value_33 <= put_Data_1_87;
          put_stuckData_4_value_34 <= put_Data_2_91;
          put_stuckData_4_value_35 <= put_Data_3_95;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        41: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        42: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        43: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2331:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        44: begin
          if (put_Found_96 >  0) begin
            put_pc <= 452;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0578:<init>|  Chip.java:0577:GONotZero|  Btree.java:2336:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        45: begin
          if (put_BtreeIndex_100 == 0) begin
            put_pc <= 47;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        46: begin
          put_pc <= 140;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        47: begin
          put_index_110 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0267:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        48: begin
          put_stuckSize_5_index_36 <= put_index_110;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_110;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_110;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_110;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        49: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        50: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        51: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        52: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        53: begin
          put_size_111 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_112 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_114 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_117 <= stuckData_stuckData_3_result_0;
          put_Key_1_118 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_121 <= stuckData_stuckData_3_result_1;
          put_Key_2_122 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_125 <= stuckData_stuckData_3_result_2;
          put_Key_3_126 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_129 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1527:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        54: begin
          if (put_size_111 < 4) begin
            put_pc <= 100;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1532:<init>|  Btree.java:1531:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        55: begin
          put_Key_0_141 <= put_Key_0_114;
          put_Data_0_144 <= put_Data_0_117;
          put_Key_1_145 <= put_Key_1_118;
          put_Data_1_148 <= put_Data_1_121;
          put_size_138 <= 2;
          put_Key_0_168 <= put_Key_2_122;
          put_Data_0_171 <= put_Data_2_125;
          put_Key_1_172 <= put_Key_3_126;
          put_Data_1_175 <= put_Data_3_129;
          put_size_165 <= 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1042:<init>|  Btree.java:1041:splitIntoTwo|  Btree.java:1549:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        56: begin
          put_root_199 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        57: begin
          put_freeNext_9_index_194 <= put_root_199;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        58: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        59: begin
          put_indexLeft_191 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        60: begin
          if (put_indexLeft_191 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_201 <= 1;
          put_isFree_202 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        61: begin
          put_freeNext_9_index_194 <= put_indexLeft_191;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_191;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_201;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_191;
          put_stuckIsFree_11_value_198 <= put_isFree_202;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        62: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        63: begin
          put_next_200 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        64: begin
          put_freeNext_10_index_195 <= put_root_199;
          put_freeNext_10_value_196 <= put_next_200;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        65: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        66: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        67: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        68: begin
          put_stuckSize_6_index_37 <= put_indexLeft_191;
          put_stuckSize_6_value_38 <= put_size_138;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_191;
          put_stuckKeys_2_value_26 <= put_Key_0_141;
          put_stuckKeys_2_value_27 <= put_Key_1_145;
          put_stuckKeys_2_value_28 <= put_Key_2_149;
          put_stuckKeys_2_value_29 <= put_Key_3_153;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_191;
          put_stuckData_4_value_32 <= put_Data_0_144;
          put_stuckData_4_value_33 <= put_Data_1_148;
          put_stuckData_4_value_34 <= put_Data_2_152;
          put_stuckData_4_value_35 <= put_Data_3_156;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        69: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        70: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        71: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1551:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        72: begin
          put_root_203 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        73: begin
          put_freeNext_9_index_194 <= put_root_203;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        74: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        75: begin
          put_indexRight_192 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        76: begin
          if (put_indexRight_192 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_205 <= 1;
          put_isFree_206 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        77: begin
          put_freeNext_9_index_194 <= put_indexRight_192;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexRight_192;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_205;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexRight_192;
          put_stuckIsFree_11_value_198 <= put_isFree_206;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        78: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        79: begin
          put_next_204 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        80: begin
          put_freeNext_10_index_195 <= put_root_203;
          put_freeNext_10_value_196 <= put_next_204;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        81: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        82: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        83: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        84: begin
          put_stuckSize_6_index_37 <= put_indexRight_192;
          put_stuckSize_6_value_38 <= put_size_165;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexRight_192;
          put_stuckKeys_2_value_26 <= put_Key_0_168;
          put_stuckKeys_2_value_27 <= put_Key_1_172;
          put_stuckKeys_2_value_28 <= put_Key_2_176;
          put_stuckKeys_2_value_29 <= put_Key_3_180;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexRight_192;
          put_stuckData_4_value_32 <= put_Data_0_171;
          put_stuckData_4_value_33 <= put_Data_1_175;
          put_stuckData_4_value_34 <= put_Data_2_179;
          put_stuckData_4_value_35 <= put_Data_3_183;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        85: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        86: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        87: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1552:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        88: begin
          case (put_size_138)
            1: begin
              put_Key_158 <= put_Key_0_141;
              put_Data_160 <= put_Data_0_144;
            end
            2: begin
              put_Key_158 <= put_Key_1_145;
              put_Data_160 <= put_Data_1_148;
            end
            3: begin
              put_Key_158 <= put_Key_2_149;
              put_Data_160 <= put_Data_2_152;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0531:<init>|  Btree.java:0530:LastElement|  Btree.java:1554:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        89: begin
          put_Key_185 <= put_Key_0_168;
          put_Data_187 <= put_Data_0_171;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0504:<init>|  Btree.java:0503:FirstElement|  Btree.java:1555:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        90: begin
          put_midKey_193 <= (put_Key_158 + put_Key_185) / 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0833:<init>|  Chip.java:0832:Average|  Btree.java:1556:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        91: begin
          put_size_111 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0395:<init>|  Btree.java:0394:Clear|  Btree.java:1557:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        92: begin
          case (put_size_111)
            0: begin
              put_Key_0_114 <= put_midKey_193;
              put_Data_0_117 <= put_indexLeft_191;
            end
            1: begin
              put_Key_1_118 <= put_midKey_193;
              put_Data_1_121 <= put_indexLeft_191;
            end
            2: begin
              put_Key_2_122 <= put_midKey_193;
              put_Data_2_125 <= put_indexLeft_191;
            end
            3: begin
              put_Key_3_126 <= put_midKey_193;
              put_Data_3_129 <= put_indexLeft_191;
            end
          endcase
          put_size_111 <= put_size_111+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0424:<init>|  Btree.java:0423:Push|  Btree.java:1558:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        93: begin
          case (put_size_111)
            0: begin
              put_Key_0_114 <= put_midKey_193;
              put_Data_0_117 <= put_indexRight_192;
            end
            1: begin
              put_Key_1_118 <= put_midKey_193;
              put_Data_1_121 <= put_indexRight_192;
            end
            2: begin
              put_Key_2_122 <= put_midKey_193;
              put_Data_2_125 <= put_indexRight_192;
            end
            3: begin
              put_Key_3_126 <= put_midKey_193;
              put_Data_3_129 <= put_indexRight_192;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0481:<init>|  Btree.java:0480:SetPastLastElement|  Btree.java:1559:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        94: begin
          put_isLeaf_112 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1560:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        95: begin
          put_stuckSize_6_index_37 <= put_index_110;
          put_stuckSize_6_value_38 <= put_size_111;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_index_110;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_112;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_110;
          put_stuckKeys_2_value_26 <= put_Key_0_114;
          put_stuckKeys_2_value_27 <= put_Key_1_118;
          put_stuckKeys_2_value_28 <= put_Key_2_122;
          put_stuckKeys_2_value_29 <= put_Key_3_126;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_110;
          put_stuckData_4_value_32 <= put_Data_0_117;
          put_stuckData_4_value_33 <= put_Data_1_121;
          put_stuckData_4_value_34 <= put_Data_2_125;
          put_stuckData_4_value_35 <= put_Data_3_129;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1561:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        96: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1561:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        97: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0329:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1561:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        98: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1561:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        99: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:1561:code|  Chip.java:0530:<init>|  Btree.java:1530:<init>|  Btree.java:1529:splitRootLeaf|  Btree.java:2340:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        100: begin
          put_BtreeIndex_100 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        101: begin
          put_index_76 <= put_BtreeIndex_100;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        102: begin
          put_stuckSize_5_index_36 <= put_index_76;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_76;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_76;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_76;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        103: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        104: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        105: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        106: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        107: begin
          put_size_77 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_78 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_80 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_83 <= stuckData_stuckData_3_result_0;
          put_Key_1_84 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_87 <= stuckData_stuckData_3_result_1;
          put_Key_2_88 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_91 <= stuckData_stuckData_3_result_2;
          put_Key_3_92 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_95 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        108: begin
          if (put_isLeaf_78 == 0) begin
            put_pc <= 115;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1395:<init>|  Btree.java:1394:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        109: begin
          put_KeyCompares_0_81 <= put_k_0 == put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 == put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 == put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 == put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0802:<init>|  Btree.java:0801:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        110: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0823:<init>|  Btree.java:0822:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        111: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0823:<init>|  Btree.java:0822:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        112: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Key_97 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Key_97 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Key_97 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Key_97 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0845:<init>|  Btree.java:0844:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        113: begin
          put_pc <= 121;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2260:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        114: begin
          put_pc <= 121;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1411:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        115: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        116: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        117: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        118: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        119: begin
          put_BtreeIndex_100 <= put_Data_99;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2264:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        120: begin
          put_pc <= 101;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2265:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        121: begin
          if (put_Found_96 == 0) begin
            put_pc <= 124;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        122: begin
          if (put_StuckIndex_101 == put_size_77) begin
            put_size_77 <= put_size_77+1;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0626:<init>|  Btree.java:0625:SetElementAt|  Btree.java:2295:Then|  Chip.java:0610:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        123: begin
          put_pc <= 135;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        124: begin
          put_notFull_208 <= put_size_77< 4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        125: begin
          if (put_notFull_208 == 0) begin
            put_pc <= 134;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        126: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        127: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        128: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        129: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        130: begin
          put_size_77 <= put_size_77+1;
          if (3 > put_StuckIndex_101) begin
            put_Key_3_92 <= put_Key_2_88;
            put_Data_3_95 <= put_Data_2_91;
          end
          if (2 > put_StuckIndex_101) begin
            put_Key_2_88 <= put_Key_1_84;
            put_Data_2_91 <= put_Data_1_87;
          end
          if (1 > put_StuckIndex_101) begin
            put_Key_1_84 <= put_Key_0_80;
            put_Data_1_87 <= put_Data_0_83;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0701:<init>|  Btree.java:0700:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        131: begin
          put_Found_96 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2305:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        132: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0592:<init>|  Chip.java:0591:COntinue|  Btree.java:2306:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        133: begin
          put_pc <= 135;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        134: begin
          put_pc <= 139;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2309:Else|  Chip.java:0620:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        135: begin
          put_stuckSize_6_index_37 <= put_index_76;
          put_stuckSize_6_value_38 <= put_size_77;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_76;
          put_stuckKeys_2_value_26 <= put_Key_0_80;
          put_stuckKeys_2_value_27 <= put_Key_1_84;
          put_stuckKeys_2_value_28 <= put_Key_2_88;
          put_stuckKeys_2_value_29 <= put_Key_3_92;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_76;
          put_stuckData_4_value_32 <= put_Data_0_83;
          put_stuckData_4_value_33 <= put_Data_1_87;
          put_stuckData_4_value_34 <= put_Data_2_91;
          put_stuckData_4_value_35 <= put_Data_3_95;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        136: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        137: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        138: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2341:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        139: begin
          put_pc <= 452;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2342:Else|  Chip.java:0620:<init>|  Btree.java:2339:<init>|  Btree.java:2338:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        140: begin
          put_index_4 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0267:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        141: begin
          put_stuckSize_5_index_36 <= put_index_4;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_4;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_4;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_4;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        142: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        143: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        144: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        145: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        146: begin
          put_size_5 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_6 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_8 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_11 <= stuckData_stuckData_3_result_0;
          put_Key_1_12 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_15 <= stuckData_stuckData_3_result_1;
          put_Key_2_16 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_19 <= stuckData_stuckData_3_result_2;
          put_Key_3_20 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_23 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:2346:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        147: begin
          put_full_107 <= put_size_5>=3 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Ge|  Btree.java:2348:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        148: begin
          if (put_full_107 == 0) begin
            put_pc <= 200;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        149: begin
          put_index_209 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0267:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        150: begin
          put_stuckSize_5_index_36 <= put_index_209;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_209;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_209;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_209;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        151: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        152: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        153: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        154: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        155: begin
          put_size_210 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_211 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_213 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_216 <= stuckData_stuckData_3_result_0;
          put_Key_1_217 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_220 <= stuckData_stuckData_3_result_1;
          put_Key_2_221 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_224 <= stuckData_stuckData_3_result_2;
          put_Key_3_225 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_228 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0268:stuckGetRoot|  Btree.java:1575:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        156: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1578:<init>|  Btree.java:1577:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        157: begin
          put_Key_0_240 <= put_Key_0_213;
          put_Data_0_243 <= put_Data_0_216;
          put_size_237 <= 1;
          put_Data_1_247 <= put_Data_1_220;
          put_Key_0_267 <= put_Key_2_221;
          put_Data_0_270 <= put_Data_2_224;
          case (put_size_210)
            0: begin
              put_size_264 <= -2;
              put_Data_1_274 <= put_Data_3_228;
            end
            1: begin
              put_size_264 <= -1;
              put_Data_1_274 <= put_Data_3_228;
            end
            2: begin
              put_size_264 <= 0;
              put_Data_1_274 <= put_Data_3_228;
            end
            3: begin
              put_size_264 <= 1;
              put_Data_1_274 <= put_Data_3_228;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1079:<init>|  Btree.java:1078:splitIntoThree|  Btree.java:1583:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        158: begin
          put_root_293 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        159: begin
          put_freeNext_9_index_194 <= put_root_293;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        160: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        161: begin
          put_indexLeft_290 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        162: begin
          if (put_indexLeft_290 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_295 <= 0;
          put_isFree_296 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        163: begin
          put_freeNext_9_index_194 <= put_indexLeft_290;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_290;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_295;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_290;
          put_stuckIsFree_11_value_198 <= put_isFree_296;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        164: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        165: begin
          put_next_294 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        166: begin
          put_freeNext_10_index_195 <= put_root_293;
          put_freeNext_10_value_196 <= put_next_294;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        167: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        168: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        169: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        170: begin
          put_stuckSize_6_index_37 <= put_indexLeft_290;
          put_stuckSize_6_value_38 <= put_size_237;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_290;
          put_stuckKeys_2_value_26 <= put_Key_0_240;
          put_stuckKeys_2_value_27 <= put_Key_1_244;
          put_stuckKeys_2_value_28 <= put_Key_2_248;
          put_stuckKeys_2_value_29 <= put_Key_3_252;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_290;
          put_stuckData_4_value_32 <= put_Data_0_243;
          put_stuckData_4_value_33 <= put_Data_1_247;
          put_stuckData_4_value_34 <= put_Data_2_251;
          put_stuckData_4_value_35 <= put_Data_3_255;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        171: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        172: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        173: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1584:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        174: begin
          put_root_297 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        175: begin
          put_freeNext_9_index_194 <= put_root_297;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        176: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        177: begin
          put_indexRight_291 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        178: begin
          if (put_indexRight_291 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_299 <= 0;
          put_isFree_300 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        179: begin
          put_freeNext_9_index_194 <= put_indexRight_291;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexRight_291;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_299;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexRight_291;
          put_stuckIsFree_11_value_198 <= put_isFree_300;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        180: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        181: begin
          put_next_298 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        182: begin
          put_freeNext_10_index_195 <= put_root_297;
          put_freeNext_10_value_196 <= put_next_298;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        183: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        184: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        185: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        186: begin
          put_stuckSize_6_index_37 <= put_indexRight_291;
          put_stuckSize_6_value_38 <= put_size_264;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexRight_291;
          put_stuckKeys_2_value_26 <= put_Key_0_267;
          put_stuckKeys_2_value_27 <= put_Key_1_271;
          put_stuckKeys_2_value_28 <= put_Key_2_275;
          put_stuckKeys_2_value_29 <= put_Key_3_279;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexRight_291;
          put_stuckData_4_value_32 <= put_Data_0_270;
          put_stuckData_4_value_33 <= put_Data_1_274;
          put_stuckData_4_value_34 <= put_Data_2_278;
          put_stuckData_4_value_35 <= put_Data_3_282;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        187: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        188: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        189: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1585:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        190: begin
          put_midKey_292 <= put_Key_1_217;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1587:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        191: begin
          put_size_210 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0395:<init>|  Btree.java:0394:Clear|  Btree.java:1588:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        192: begin
          case (put_size_210)
            0: begin
              put_Key_0_213 <= put_midKey_292;
              put_Data_0_216 <= put_indexLeft_290;
            end
            1: begin
              put_Key_1_217 <= put_midKey_292;
              put_Data_1_220 <= put_indexLeft_290;
            end
            2: begin
              put_Key_2_221 <= put_midKey_292;
              put_Data_2_224 <= put_indexLeft_290;
            end
            3: begin
              put_Key_3_225 <= put_midKey_292;
              put_Data_3_228 <= put_indexLeft_290;
            end
          endcase
          put_size_210 <= put_size_210+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0424:<init>|  Btree.java:0423:Push|  Btree.java:1589:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        193: begin
          case (put_size_210)
            0: begin
              put_Key_0_213 <= put_midKey_292;
              put_Data_0_216 <= put_indexRight_291;
            end
            1: begin
              put_Key_1_217 <= put_midKey_292;
              put_Data_1_220 <= put_indexRight_291;
            end
            2: begin
              put_Key_2_221 <= put_midKey_292;
              put_Data_2_224 <= put_indexRight_291;
            end
            3: begin
              put_Key_3_225 <= put_midKey_292;
              put_Data_3_228 <= put_indexRight_291;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0481:<init>|  Btree.java:0480:SetPastLastElement|  Btree.java:1590:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        194: begin
          put_stuckSize_6_index_37 <= put_index_209;
          put_stuckSize_6_value_38 <= put_size_210;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_209;
          put_stuckKeys_2_value_26 <= put_Key_0_213;
          put_stuckKeys_2_value_27 <= put_Key_1_217;
          put_stuckKeys_2_value_28 <= put_Key_2_221;
          put_stuckKeys_2_value_29 <= put_Key_3_225;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_209;
          put_stuckData_4_value_32 <= put_Data_0_216;
          put_stuckData_4_value_33 <= put_Data_1_220;
          put_stuckData_4_value_34 <= put_Data_2_224;
          put_stuckData_4_value_35 <= put_Data_3_228;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1591:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        195: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1591:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        196: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1591:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        197: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1591:splitRootBranch|  Btree.java:2352:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        198: begin
          put_pc <= 44;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2353:Then|  Chip.java:0610:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        199: begin
          put_pc <= 200;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2351:<init>|  Btree.java:2350:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        200: begin
          put_parent_104 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2357:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        201: begin
          put_index_4 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        202: begin
          put_stuckSize_5_index_36 <= put_index_4;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_4;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_4;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_4;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        203: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        204: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        205: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        206: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        207: begin
          put_size_5 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_6 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_8 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_11 <= stuckData_stuckData_3_result_0;
          put_Key_1_12 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_15 <= stuckData_stuckData_3_result_1;
          put_Key_2_16 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_19 <= stuckData_stuckData_3_result_2;
          put_Key_3_20 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_23 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2362:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        208: begin
          put_KeyCompares_0_9 <= put_k_0 <= put_Key_0_8 && 0 < put_size_5;
          put_KeyCollapse_0_10 <= 0;
          put_KeyCompares_1_13 <= put_k_0 >  put_Key_0_8 && put_k_0 <= put_Key_1_12 && 1 < put_size_5;
          put_KeyCollapse_1_14 <= 1;
          put_KeyCompares_2_17 <= put_k_0 >  put_Key_1_12 && put_k_0 <= put_Key_2_16 && 2 < put_size_5;
          put_KeyCollapse_2_18 <= 2;
          put_KeyCompares_3_21 <= put_k_0 >  put_Key_2_16 && put_k_0 <= put_Key_3_20 && 3 < put_size_5;
          put_KeyCollapse_3_22 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2363:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        209: begin
          if (put_KeyCompares_1_13) begin
            put_KeyCompares_0_9 <= 1;
            put_KeyCollapse_0_10 <= put_KeyCollapse_1_14;
          end
          if (put_KeyCompares_3_21) begin
            put_KeyCompares_2_17 <= 1;
            put_KeyCollapse_2_18 <= put_KeyCollapse_3_22;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2363:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        210: begin
          if (put_KeyCompares_2_17) begin
            put_KeyCompares_0_9 <= 1;
            put_KeyCollapse_0_10 <= put_KeyCollapse_2_18;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2363:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        211: begin
          if (put_KeyCompares_0_9) begin
            put_Found_42 <= 1;
            case (put_KeyCollapse_0_10)
              0: begin
                put_StuckIndex_47 <= 0;
                put_FoundKey_44 <= put_Key_0_8;
                put_Data_45 <= put_Data_0_11;
              end
              1: begin
                put_StuckIndex_47 <= 1;
                put_FoundKey_44 <= put_Key_1_12;
                put_Data_45 <= put_Data_1_15;
              end
              2: begin
                put_StuckIndex_47 <= 2;
                put_FoundKey_44 <= put_Key_2_16;
                put_Data_45 <= put_Data_2_19;
              end
              3: begin
                put_StuckIndex_47 <= 3;
                put_FoundKey_44 <= put_Key_3_20;
                put_Data_45 <= put_Data_3_23;
              end
            endcase
          end
          else begin
            put_Found_42 <= 0;
            case (put_size_5)
              0: begin
                put_StuckIndex_47 <= 0;
                put_Data_45 <= put_Data_0_11;
              end
              1: begin
                put_StuckIndex_47 <= 1;
                put_Data_45 <= put_Data_1_15;
              end
              2: begin
                put_StuckIndex_47 <= 2;
                put_Data_45 <= put_Data_2_19;
              end
              3: begin
                put_StuckIndex_47 <= 3;
                put_Data_45 <= put_Data_3_23;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2363:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        212: begin
          put_child_103 <= put_Data_45;
          put_childInparent_105 <= put_StuckIndex_47;
          put_found_106 <= put_Found_42;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2365:<init>|  Btree.java:2364:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        213: begin
          put_index_49 <= put_child_103;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        214: begin
          put_stuckSize_5_index_36 <= put_index_49;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_49;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_49;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_49;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        215: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        216: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        217: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        218: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        219: begin
          put_size_50 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_51 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_53 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_56 <= stuckData_stuckData_3_result_0;
          put_Key_1_57 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_60 <= stuckData_stuckData_3_result_1;
          put_Key_2_61 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_64 <= stuckData_stuckData_3_result_2;
          put_Key_3_65 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_68 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2373:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        220: begin
          if (put_isLeaf_51 == 0) begin
            put_pc <= 359;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1395:<init>|  Btree.java:1394:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        221: begin
          put_full_107 <= put_size_50>=4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Ge|  Btree.java:2377:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        222: begin
          if (put_full_107 == 0) begin
            put_pc <= 318;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        223: begin
          if (put_found_106 == 0) begin
            put_pc <= 270;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        224: begin
          put_index_301 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        225: begin
          put_stuckSize_5_index_36 <= put_index_301;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_301;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_301;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_301;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        226: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        227: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        228: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        229: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        230: begin
          put_size_302 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_303 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_305 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_308 <= stuckData_stuckData_3_result_0;
          put_Key_1_309 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_312 <= stuckData_stuckData_3_result_1;
          put_Key_2_313 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_316 <= stuckData_stuckData_3_result_2;
          put_Key_3_317 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_320 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1607:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        231: begin
          case (put_childInparent_105)
            0: begin
              put_childKey_409 <= put_Key_0_305;
              put_childData_410 <= put_Data_0_308;
            end
            1: begin
              put_childKey_409 <= put_Key_1_309;
              put_childData_410 <= put_Data_1_312;
            end
            2: begin
              put_childKey_409 <= put_Key_2_313;
              put_childData_410 <= put_Data_2_316;
            end
            3: begin
              put_childKey_409 <= put_Key_3_317;
              put_childData_410 <= put_Data_3_320;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1610:<init>|  Btree.java:1609:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        232: begin
          put_index_328 <= put_childData_410;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        233: begin
          put_stuckSize_5_index_36 <= put_index_328;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_328;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_328;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_328;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        234: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        235: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        236: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        237: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        238: begin
          put_size_329 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_330 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_332 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_335 <= stuckData_stuckData_3_result_0;
          put_Key_1_336 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_339 <= stuckData_stuckData_3_result_1;
          put_Key_2_340 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_343 <= stuckData_stuckData_3_result_2;
          put_Key_3_344 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_347 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1623:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        239: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1626:<init>|  Btree.java:1625:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        240: begin
          put_Key_0_359 <= put_Key_0_332;
          put_Data_0_362 <= put_Data_0_335;
          put_Key_1_363 <= put_Key_1_336;
          put_Data_1_366 <= put_Data_1_339;
          put_size_356 <= 2;
          put_Key_0_332 <= put_Key_2_340;
          put_Data_0_335 <= put_Data_2_343;
          put_Key_1_336 <= put_Key_3_344;
          put_Data_1_339 <= put_Data_3_347;
          put_size_329 <= 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1125:<init>|  Btree.java:1124:splitLow|  Btree.java:1634:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        241: begin
          put_root_414 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        242: begin
          put_freeNext_9_index_194 <= put_root_414;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        243: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        244: begin
          put_indexLeft_411 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        245: begin
          if (put_indexLeft_411 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_416 <= 1;
          put_isFree_417 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        246: begin
          put_freeNext_9_index_194 <= put_indexLeft_411;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_411;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_416;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_411;
          put_stuckIsFree_11_value_198 <= put_isFree_417;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        247: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        248: begin
          put_next_415 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        249: begin
          put_freeNext_10_index_195 <= put_root_414;
          put_freeNext_10_value_196 <= put_next_415;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        250: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        251: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        252: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        253: begin
          put_stuckSize_6_index_37 <= put_childData_410;
          put_stuckSize_6_value_38 <= put_size_329;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childData_410;
          put_stuckKeys_2_value_26 <= put_Key_0_332;
          put_stuckKeys_2_value_27 <= put_Key_1_336;
          put_stuckKeys_2_value_28 <= put_Key_2_340;
          put_stuckKeys_2_value_29 <= put_Key_3_344;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childData_410;
          put_stuckData_4_value_32 <= put_Data_0_335;
          put_stuckData_4_value_33 <= put_Data_1_339;
          put_stuckData_4_value_34 <= put_Data_2_343;
          put_stuckData_4_value_35 <= put_Data_3_347;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        254: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        255: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        256: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1635:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        257: begin
          put_stuckSize_6_index_37 <= put_indexLeft_411;
          put_stuckSize_6_value_38 <= put_size_356;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_411;
          put_stuckKeys_2_value_26 <= put_Key_0_359;
          put_stuckKeys_2_value_27 <= put_Key_1_363;
          put_stuckKeys_2_value_28 <= put_Key_2_367;
          put_stuckKeys_2_value_29 <= put_Key_3_371;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_411;
          put_stuckData_4_value_32 <= put_Data_0_362;
          put_stuckData_4_value_33 <= put_Data_1_366;
          put_stuckData_4_value_34 <= put_Data_2_370;
          put_stuckData_4_value_35 <= put_Data_3_374;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1636:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        258: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1636:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        259: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1636:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        260: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1636:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        261: begin
          case (put_size_356)
            1: begin
              put_Key_376 <= put_Key_0_359;
              put_Data_378 <= put_Data_0_362;
            end
            2: begin
              put_Key_376 <= put_Key_1_363;
              put_Data_378 <= put_Data_1_366;
            end
            3: begin
              put_Key_376 <= put_Key_2_367;
              put_Data_378 <= put_Data_2_370;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0531:<init>|  Btree.java:0530:LastElement|  Btree.java:1638:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        262: begin
          put_Key_349 <= put_Key_0_332;
          put_Data_351 <= put_Data_0_335;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0504:<init>|  Btree.java:0503:FirstElement|  Btree.java:1639:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        263: begin
          put_midKey_413 <= (put_Key_376 + put_Key_349) / 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0833:<init>|  Chip.java:0832:Average|  Btree.java:1640:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        264: begin
          put_size_302 <= put_size_302+1;
          if (3 > put_childInparent_105) begin
            put_Key_3_317 <= put_Key_2_313;
            put_Data_3_320 <= put_Data_2_316;
          end
          if (2 > put_childInparent_105) begin
            put_Key_2_313 <= put_Key_1_309;
            put_Data_2_316 <= put_Data_1_312;
          end
          if (1 > put_childInparent_105) begin
            put_Key_1_309 <= put_Key_0_305;
            put_Data_1_312 <= put_Data_0_308;
          end
          case (put_childInparent_105)
            0: begin
              put_Key_0_305 <= put_midKey_413;
              put_Data_0_308 <= put_indexLeft_411;
            end
            1: begin
              put_Key_1_309 <= put_midKey_413;
              put_Data_1_312 <= put_indexLeft_411;
            end
            2: begin
              put_Key_2_313 <= put_midKey_413;
              put_Data_2_316 <= put_indexLeft_411;
            end
            3: begin
              put_Key_3_317 <= put_midKey_413;
              put_Data_3_320 <= put_indexLeft_411;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0701:<init>|  Btree.java:0700:InsertElementAt|  Btree.java:1641:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        265: begin
          put_stuckSize_6_index_37 <= put_index_301;
          put_stuckSize_6_value_38 <= put_size_302;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_301;
          put_stuckKeys_2_value_26 <= put_Key_0_305;
          put_stuckKeys_2_value_27 <= put_Key_1_309;
          put_stuckKeys_2_value_28 <= put_Key_2_313;
          put_stuckKeys_2_value_29 <= put_Key_3_317;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_301;
          put_stuckData_4_value_32 <= put_Data_0_308;
          put_stuckData_4_value_33 <= put_Data_1_312;
          put_stuckData_4_value_34 <= put_Data_2_316;
          put_stuckData_4_value_35 <= put_Data_3_320;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1642:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        266: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1642:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        267: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1642:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        268: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1642:splitLeafNotTop|  Btree.java:2383:Then|  Chip.java:0610:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        269: begin
          put_pc <= 317;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        270: begin
          put_index_418 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        271: begin
          put_stuckSize_5_index_36 <= put_index_418;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_418;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_418;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_418;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        272: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        273: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        274: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        275: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        276: begin
          put_size_419 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_420 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_422 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_425 <= stuckData_stuckData_3_result_0;
          put_Key_1_426 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_429 <= stuckData_stuckData_3_result_1;
          put_Key_2_430 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_433 <= stuckData_stuckData_3_result_2;
          put_Key_3_434 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_437 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1654:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        277: begin
          case (put_size_419)
            0: begin
              put_Key_439 <= put_Key_0_422;
              put_Data_441 <= put_Data_0_425;
            end
            1: begin
              put_Key_439 <= put_Key_1_426;
              put_Data_441 <= put_Data_1_429;
            end
            2: begin
              put_Key_439 <= put_Key_2_430;
              put_Data_441 <= put_Data_2_433;
            end
            3: begin
              put_Key_439 <= put_Key_3_434;
              put_Data_441 <= put_Data_3_437;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0558:<init>|  Btree.java:0557:PastLastElement|  Btree.java:1655:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        278: begin
          put_childIndex_499 <= put_Data_441;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1656:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        279: begin
          put_index_445 <= put_childIndex_499;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        280: begin
          put_stuckSize_5_index_36 <= put_index_445;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_445;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_445;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_445;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        281: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        282: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        283: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        284: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        285: begin
          put_size_446 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_447 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_449 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_452 <= stuckData_stuckData_3_result_0;
          put_Key_1_453 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_456 <= stuckData_stuckData_3_result_1;
          put_Key_2_457 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_460 <= stuckData_stuckData_3_result_2;
          put_Key_3_461 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_464 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1657:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        286: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1660:<init>|  Btree.java:1659:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        287: begin
          put_Key_0_476 <= put_Key_0_449;
          put_Data_0_479 <= put_Data_0_452;
          put_Key_1_480 <= put_Key_1_453;
          put_Data_1_483 <= put_Data_1_456;
          put_size_473 <= 2;
          put_Key_0_449 <= put_Key_2_457;
          put_Data_0_452 <= put_Data_2_460;
          put_Key_1_453 <= put_Key_3_461;
          put_Data_1_456 <= put_Data_3_464;
          put_size_446 <= 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1125:<init>|  Btree.java:1124:splitLow|  Btree.java:1669:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        288: begin
          put_root_502 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        289: begin
          put_freeNext_9_index_194 <= put_root_502;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        290: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        291: begin
          put_leftIndex_500 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        292: begin
          if (put_leftIndex_500 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_504 <= 1;
          put_isFree_505 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        293: begin
          put_freeNext_9_index_194 <= put_leftIndex_500;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_leftIndex_500;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_504;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_leftIndex_500;
          put_stuckIsFree_11_value_198 <= put_isFree_505;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        294: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        295: begin
          put_next_503 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        296: begin
          put_freeNext_10_index_195 <= put_root_502;
          put_freeNext_10_value_196 <= put_next_503;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        297: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        298: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        299: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0151:allocateLeaf|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        300: begin
          put_stuckSize_6_index_37 <= put_leftIndex_500;
          put_stuckSize_6_value_38 <= put_size_473;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_leftIndex_500;
          put_stuckKeys_2_value_26 <= put_Key_0_476;
          put_stuckKeys_2_value_27 <= put_Key_1_480;
          put_stuckKeys_2_value_28 <= put_Key_2_484;
          put_stuckKeys_2_value_29 <= put_Key_3_488;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_leftIndex_500;
          put_stuckData_4_value_32 <= put_Data_0_479;
          put_stuckData_4_value_33 <= put_Data_1_483;
          put_stuckData_4_value_34 <= put_Data_2_487;
          put_stuckData_4_value_35 <= put_Data_3_491;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        301: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        302: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        303: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        304: begin
          put_stuckSize_6_index_37 <= put_childIndex_499;
          put_stuckSize_6_value_38 <= put_size_446;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childIndex_499;
          put_stuckKeys_2_value_26 <= put_Key_0_449;
          put_stuckKeys_2_value_27 <= put_Key_1_453;
          put_stuckKeys_2_value_28 <= put_Key_2_457;
          put_stuckKeys_2_value_29 <= put_Key_3_461;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childIndex_499;
          put_stuckData_4_value_32 <= put_Data_0_452;
          put_stuckData_4_value_33 <= put_Data_1_456;
          put_stuckData_4_value_34 <= put_Data_2_460;
          put_stuckData_4_value_35 <= put_Data_3_464;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        305: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        306: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        307: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1670:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        308: begin
          case (put_size_473)
            1: begin
              put_Key_493 <= put_Key_0_476;
              put_Data_495 <= put_Data_0_479;
            end
            2: begin
              put_Key_493 <= put_Key_1_480;
              put_Data_495 <= put_Data_1_483;
            end
            3: begin
              put_Key_493 <= put_Key_2_484;
              put_Data_495 <= put_Data_2_487;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0531:<init>|  Btree.java:0530:LastElement|  Btree.java:1672:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        309: begin
          put_Key_466 <= put_Key_0_449;
          put_Data_468 <= put_Data_0_452;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0504:<init>|  Btree.java:0503:FirstElement|  Btree.java:1673:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        310: begin
          put_midKey_501 <= (put_Key_493 + put_Key_466) / 2;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0833:<init>|  Chip.java:0832:Average|  Btree.java:1674:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        311: begin
          case (put_size_419)
            0: begin
              put_Key_0_422 <= put_midKey_501;
              put_Data_0_425 <= put_leftIndex_500;
            end
            1: begin
              put_Key_1_426 <= put_midKey_501;
              put_Data_1_429 <= put_leftIndex_500;
            end
            2: begin
              put_Key_2_430 <= put_midKey_501;
              put_Data_2_433 <= put_leftIndex_500;
            end
            3: begin
              put_Key_3_434 <= put_midKey_501;
              put_Data_3_437 <= put_leftIndex_500;
            end
          endcase
          put_size_419 <= put_size_419+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0424:<init>|  Btree.java:0423:Push|  Btree.java:1675:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        312: begin
          case (put_size_419)
            0: begin
              put_Key_0_422 <= put_midKey_501;
              put_Data_0_425 <= put_childIndex_499;
            end
            1: begin
              put_Key_1_426 <= put_midKey_501;
              put_Data_1_429 <= put_childIndex_499;
            end
            2: begin
              put_Key_2_430 <= put_midKey_501;
              put_Data_2_433 <= put_childIndex_499;
            end
            3: begin
              put_Key_3_434 <= put_midKey_501;
              put_Data_3_437 <= put_childIndex_499;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0481:<init>|  Btree.java:0480:SetPastLastElement|  Btree.java:1676:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        313: begin
          put_stuckSize_6_index_37 <= put_index_418;
          put_stuckSize_6_value_38 <= put_size_419;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_418;
          put_stuckKeys_2_value_26 <= put_Key_0_422;
          put_stuckKeys_2_value_27 <= put_Key_1_426;
          put_stuckKeys_2_value_28 <= put_Key_2_430;
          put_stuckKeys_2_value_29 <= put_Key_3_434;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_418;
          put_stuckData_4_value_32 <= put_Data_0_425;
          put_stuckData_4_value_33 <= put_Data_1_429;
          put_stuckData_4_value_34 <= put_Data_2_433;
          put_stuckData_4_value_35 <= put_Data_3_437;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        314: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        315: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        316: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1677:splitLeafAtTop|  Btree.java:2386:Else|  Chip.java:0620:<init>|  Btree.java:2382:<init>|  Btree.java:2381:Then|  Chip.java:0610:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        317: begin
          put_pc <= 318;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2380:<init>|  Btree.java:2379:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        318: begin
          put_BtreeIndex_100 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2252:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        319: begin
          put_index_76 <= put_BtreeIndex_100;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        320: begin
          put_stuckSize_5_index_36 <= put_index_76;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_76;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_76;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_76;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        321: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        322: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        323: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        324: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        325: begin
          put_size_77 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_78 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_80 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_83 <= stuckData_stuckData_3_result_0;
          put_Key_1_84 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_87 <= stuckData_stuckData_3_result_1;
          put_Key_2_88 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_91 <= stuckData_stuckData_3_result_2;
          put_Key_3_92 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_95 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:2256:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        326: begin
          if (put_isLeaf_78 == 0) begin
            put_pc <= 333;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1395:<init>|  Btree.java:1394:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        327: begin
          put_KeyCompares_0_81 <= put_k_0 == put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 == put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 == put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 == put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0802:<init>|  Btree.java:0801:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        328: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0823:<init>|  Btree.java:0822:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        329: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0823:<init>|  Btree.java:0822:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        330: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Key_97 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Key_97 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Key_97 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Key_97 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0845:<init>|  Btree.java:0844:search_eq_parallel|  Btree.java:2259:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        331: begin
          put_pc <= 339;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2260:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        332: begin
          put_pc <= 339;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1411:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        333: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        334: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        335: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        336: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2263:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        337: begin
          put_BtreeIndex_100 <= put_Data_99;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2264:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        338: begin
          put_pc <= 319;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2265:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2258:<init>|  Btree.java:2257:code|  Chip.java:0530:<init>|  Btree.java:2255:<init>|  Btree.java:2254:findSearch|  Btree.java:2291:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        339: begin
          if (put_Found_96 == 0) begin
            put_pc <= 342;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        340: begin
          if (put_StuckIndex_101 == put_size_77) begin
            put_size_77 <= put_size_77+1;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0626:<init>|  Btree.java:0625:SetElementAt|  Btree.java:2295:Then|  Chip.java:0610:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        341: begin
          put_pc <= 353;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        342: begin
          put_notFull_507 <= put_size_77< 4 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:2299:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        343: begin
          if (put_notFull_507 == 0) begin
            put_pc <= 352;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        344: begin
          put_KeyCompares_0_81 <= put_k_0 <= put_Key_0_80 && 0 < put_size_77;
          put_KeyCollapse_0_82 <= 0;
          put_KeyCompares_1_85 <= put_k_0 >  put_Key_0_80 && put_k_0 <= put_Key_1_84 && 1 < put_size_77;
          put_KeyCollapse_1_86 <= 1;
          put_KeyCompares_2_89 <= put_k_0 >  put_Key_1_84 && put_k_0 <= put_Key_2_88 && 2 < put_size_77;
          put_KeyCollapse_2_90 <= 2;
          put_KeyCompares_3_93 <= put_k_0 >  put_Key_2_88 && put_k_0 <= put_Key_3_92 && 3 < put_size_77;
          put_KeyCollapse_3_94 <= 3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0938:<init>|  Btree.java:0937:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        345: begin
          if (put_KeyCompares_1_85) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_1_86;
          end
          if (put_KeyCompares_3_93) begin
            put_KeyCompares_2_89 <= 1;
            put_KeyCollapse_2_90 <= put_KeyCollapse_3_94;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        346: begin
          if (put_KeyCompares_2_89) begin
            put_KeyCompares_0_81 <= 1;
            put_KeyCollapse_0_82 <= put_KeyCollapse_2_90;
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0974:<init>|  Btree.java:0973:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        347: begin
          if (put_KeyCompares_0_81) begin
            put_Found_96 <= 1;
            case (put_KeyCollapse_0_82)
              0: begin
                put_StuckIndex_101 <= 0;
                put_FoundKey_98 <= put_Key_0_80;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_FoundKey_98 <= put_Key_1_84;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_FoundKey_98 <= put_Key_2_88;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_FoundKey_98 <= put_Key_3_92;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          else begin
            put_Found_96 <= 0;
            case (put_size_77)
              0: begin
                put_StuckIndex_101 <= 0;
                put_Data_99 <= put_Data_0_83;
              end
              1: begin
                put_StuckIndex_101 <= 1;
                put_Data_99 <= put_Data_1_87;
              end
              2: begin
                put_StuckIndex_101 <= 2;
                put_Data_99 <= put_Data_2_91;
              end
              3: begin
                put_StuckIndex_101 <= 3;
                put_Data_99 <= put_Data_3_95;
              end
            endcase
          end
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0996:<init>|  Btree.java:0995:search_le_parallel|  Btree.java:2303:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        348: begin
          put_size_77 <= put_size_77+1;
          if (3 > put_StuckIndex_101) begin
            put_Key_3_92 <= put_Key_2_88;
            put_Data_3_95 <= put_Data_2_91;
          end
          if (2 > put_StuckIndex_101) begin
            put_Key_2_88 <= put_Key_1_84;
            put_Data_2_91 <= put_Data_1_87;
          end
          if (1 > put_StuckIndex_101) begin
            put_Key_1_84 <= put_Key_0_80;
            put_Data_1_87 <= put_Data_0_83;
          end
          case (put_StuckIndex_101)
            0: begin
              put_Key_0_80 <= put_k_0;
              put_Data_0_83 <= put_d_1;
            end
            1: begin
              put_Key_1_84 <= put_k_0;
              put_Data_1_87 <= put_d_1;
            end
            2: begin
              put_Key_2_88 <= put_k_0;
              put_Data_2_91 <= put_d_1;
            end
            3: begin
              put_Key_3_92 <= put_k_0;
              put_Data_3_95 <= put_d_1;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0701:<init>|  Btree.java:0700:InsertElementAt|  Btree.java:2304:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        349: begin
          put_Found_96 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0799:<init>|  Chip.java:0798:One|  Btree.java:2305:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        350: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0592:<init>|  Chip.java:0591:COntinue|  Btree.java:2306:Then|  Chip.java:0610:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        351: begin
          put_pc <= 353;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        352: begin
          put_pc <= 357;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2309:Else|  Chip.java:0620:<init>|  Btree.java:2302:<init>|  Btree.java:2301:Else|  Chip.java:0620:<init>|  Btree.java:2294:<init>|  Btree.java:2293:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        353: begin
          put_stuckSize_6_index_37 <= put_index_76;
          put_stuckSize_6_value_38 <= put_size_77;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_76;
          put_stuckKeys_2_value_26 <= put_Key_0_80;
          put_stuckKeys_2_value_27 <= put_Key_1_84;
          put_stuckKeys_2_value_28 <= put_Key_2_88;
          put_stuckKeys_2_value_29 <= put_Key_3_92;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_76;
          put_stuckData_4_value_32 <= put_Data_0_83;
          put_stuckData_4_value_33 <= put_Data_1_87;
          put_stuckData_4_value_34 <= put_Data_2_91;
          put_stuckData_4_value_35 <= put_Data_3_95;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        354: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        355: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        356: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0337:stuckPut|  Btree.java:2314:code|  Chip.java:0530:<init>|  Btree.java:2290:<init>|  Btree.java:2289:findAndInsert|  Btree.java:2391:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        357: begin
          put_pc <= 452;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2392:Leaf|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        358: begin
          put_pc <= 452;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1411:code|  Chip.java:0530:<init>|  Btree.java:1392:<init>|  Btree.java:1391:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        359: begin
          put_full_107 <= put_size_50>=3 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0784:<init>|  Chip.java:0784:Ge|  Btree.java:2396:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        360: begin
          if (put_full_107 == 0) begin
            put_pc <= 450;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        361: begin
          if (put_found_106 == 0) begin
            put_pc <= 405;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        362: begin
          put_index_508 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        363: begin
          put_stuckSize_5_index_36 <= put_index_508;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_508;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_508;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_508;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        364: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        365: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        366: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        367: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        368: begin
          put_size_509 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_510 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_512 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_515 <= stuckData_stuckData_3_result_0;
          put_Key_1_516 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_519 <= stuckData_stuckData_3_result_1;
          put_Key_2_520 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_523 <= stuckData_stuckData_3_result_2;
          put_Key_3_524 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_527 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1693:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        369: begin
          case (put_childInparent_105)
            0: begin
              put_childKey_616 <= put_Key_0_512;
              put_childData_617 <= put_Data_0_515;
            end
            1: begin
              put_childKey_616 <= put_Key_1_516;
              put_childData_617 <= put_Data_1_519;
            end
            2: begin
              put_childKey_616 <= put_Key_2_520;
              put_childData_617 <= put_Data_2_523;
            end
            3: begin
              put_childKey_616 <= put_Key_3_524;
              put_childData_617 <= put_Data_3_527;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1695:<init>|  Btree.java:1694:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        370: begin
          put_index_535 <= put_childData_617;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        371: begin
          put_stuckSize_5_index_36 <= put_index_535;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_535;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_535;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_535;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        372: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        373: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        374: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        375: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        376: begin
          put_size_536 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_537 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_539 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_542 <= stuckData_stuckData_3_result_0;
          put_Key_1_543 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_546 <= stuckData_stuckData_3_result_1;
          put_Key_2_547 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_550 <= stuckData_stuckData_3_result_2;
          put_Key_3_551 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_554 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1708:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        377: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1711:<init>|  Btree.java:1710:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        378: begin
          put_Key_0_566 <= put_Key_0_539;
          put_Data_0_569 <= put_Data_0_542;
          put_size_563 <= 1;
          put_Data_1_573 <= put_Data_1_546;
          put_childKey_616 <= put_Key_1_543;
          put_Key_0_539 <= put_Key_2_547;
          put_Data_0_542 <= put_Data_2_550;
          put_Key_1_543 <= put_Key_3_551;
          put_Data_1_546 <= put_Data_3_554;
          put_size_536 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1166:<init>|  Btree.java:1165:splitLowButOne|  Btree.java:1720:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        379: begin
          put_root_621 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        380: begin
          put_freeNext_9_index_194 <= put_root_621;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        381: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        382: begin
          put_indexLeft_618 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        383: begin
          if (put_indexLeft_618 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_623 <= 0;
          put_isFree_624 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        384: begin
          put_freeNext_9_index_194 <= put_indexLeft_618;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_618;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_623;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_618;
          put_stuckIsFree_11_value_198 <= put_isFree_624;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        385: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        386: begin
          put_next_622 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        387: begin
          put_freeNext_10_index_195 <= put_root_621;
          put_freeNext_10_value_196 <= put_next_622;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        388: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        389: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        390: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        391: begin
          put_stuckSize_6_index_37 <= put_indexLeft_618;
          put_stuckSize_6_value_38 <= put_size_563;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_618;
          put_stuckKeys_2_value_26 <= put_Key_0_566;
          put_stuckKeys_2_value_27 <= put_Key_1_570;
          put_stuckKeys_2_value_28 <= put_Key_2_574;
          put_stuckKeys_2_value_29 <= put_Key_3_578;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_618;
          put_stuckData_4_value_32 <= put_Data_0_569;
          put_stuckData_4_value_33 <= put_Data_1_573;
          put_stuckData_4_value_34 <= put_Data_2_577;
          put_stuckData_4_value_35 <= put_Data_3_581;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        392: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        393: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        394: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1721:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        395: begin
          put_stuckSize_6_index_37 <= put_childData_617;
          put_stuckSize_6_value_38 <= put_size_536;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childData_617;
          put_stuckKeys_2_value_26 <= put_Key_0_539;
          put_stuckKeys_2_value_27 <= put_Key_1_543;
          put_stuckKeys_2_value_28 <= put_Key_2_547;
          put_stuckKeys_2_value_29 <= put_Key_3_551;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childData_617;
          put_stuckData_4_value_32 <= put_Data_0_542;
          put_stuckData_4_value_33 <= put_Data_1_546;
          put_stuckData_4_value_34 <= put_Data_2_550;
          put_stuckData_4_value_35 <= put_Data_3_554;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1722:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        396: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1722:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        397: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1722:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        398: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1722:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        399: begin
          put_size_509 <= put_size_509+1;
          if (3 > put_childInparent_105) begin
            put_Key_3_524 <= put_Key_2_520;
            put_Data_3_527 <= put_Data_2_523;
          end
          if (2 > put_childInparent_105) begin
            put_Key_2_520 <= put_Key_1_516;
            put_Data_2_523 <= put_Data_1_519;
          end
          if (1 > put_childInparent_105) begin
            put_Key_1_516 <= put_Key_0_512;
            put_Data_1_519 <= put_Data_0_515;
          end
          case (put_childInparent_105)
            0: begin
              put_Key_0_512 <= put_childKey_616;
              put_Data_0_515 <= put_indexLeft_618;
            end
            1: begin
              put_Key_1_516 <= put_childKey_616;
              put_Data_1_519 <= put_indexLeft_618;
            end
            2: begin
              put_Key_2_520 <= put_childKey_616;
              put_Data_2_523 <= put_indexLeft_618;
            end
            3: begin
              put_Key_3_524 <= put_childKey_616;
              put_Data_3_527 <= put_indexLeft_618;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0701:<init>|  Btree.java:0700:InsertElementAt|  Btree.java:1724:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        400: begin
          put_stuckSize_6_index_37 <= put_index_508;
          put_stuckSize_6_value_38 <= put_size_509;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_508;
          put_stuckKeys_2_value_26 <= put_Key_0_512;
          put_stuckKeys_2_value_27 <= put_Key_1_516;
          put_stuckKeys_2_value_28 <= put_Key_2_520;
          put_stuckKeys_2_value_29 <= put_Key_3_524;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_508;
          put_stuckData_4_value_32 <= put_Data_0_515;
          put_stuckData_4_value_33 <= put_Data_1_519;
          put_stuckData_4_value_34 <= put_Data_2_523;
          put_stuckData_4_value_35 <= put_Data_3_527;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1725:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        401: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1725:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        402: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1725:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        403: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1725:splitBranchNotTop|  Btree.java:2402:Then|  Chip.java:0610:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        404: begin
          put_pc <= 449;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        405: begin
          put_index_625 <= put_parent_104;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        406: begin
          put_stuckSize_5_index_36 <= put_index_625;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_625;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_625;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_625;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        407: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        408: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        409: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        410: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        411: begin
          put_size_626 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_627 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_629 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_632 <= stuckData_stuckData_3_result_0;
          put_Key_1_633 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_636 <= stuckData_stuckData_3_result_1;
          put_Key_2_637 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_640 <= stuckData_stuckData_3_result_2;
          put_Key_3_641 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_644 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1740:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        412: begin
          case (put_size_626)
            0: begin
              put_Key_646 <= put_Key_0_629;
              put_Data_648 <= put_Data_0_632;
            end
            1: begin
              put_Key_646 <= put_Key_1_633;
              put_Data_648 <= put_Data_1_636;
            end
            2: begin
              put_Key_646 <= put_Key_2_637;
              put_Data_648 <= put_Data_2_640;
            end
            3: begin
              put_Key_646 <= put_Key_3_641;
              put_Data_648 <= put_Data_3_644;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0558:<init>|  Btree.java:0557:PastLastElement|  Btree.java:1742:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        413: begin
          put_childData_734 <= put_Data_648;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:1743:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        414: begin
          put_index_652 <= put_childData_734;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0262:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        415: begin
          put_stuckSize_5_index_36 <= put_index_652;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          put_stuckIsLeaf_7_index_39 <= put_index_652;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          put_stuckKeys_1_index_24 <= put_index_652;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          put_stuckData_3_index_30 <= put_index_652;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0273:<init>|  Btree.java:0272:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        416: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        417: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0287:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        418: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        419: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0290:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        420: begin
          put_size_653 <= stuckSize_stuckSize_5_result_0;
          put_isLeaf_654 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          put_Key_0_656 <= stuckKeys_stuckKeys_1_result_0;
          put_Data_0_659 <= stuckData_stuckData_3_result_0;
          put_Key_1_660 <= stuckKeys_stuckKeys_1_result_1;
          put_Data_1_663 <= stuckData_stuckData_3_result_1;
          put_Key_2_664 <= stuckKeys_stuckKeys_1_result_2;
          put_Data_2_667 <= stuckData_stuckData_3_result_2;
          put_Key_3_668 <= stuckKeys_stuckKeys_1_result_3;
          put_Data_3_671 <= stuckData_stuckData_3_result_3;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0293:<init>|  Btree.java:0292:stuckGet|  Btree.java:0263:stuckGet|  Btree.java:1744:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        421: begin
          
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1747:<init>|  Btree.java:1746:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        422: begin
          put_Key_0_683 <= put_Key_0_656;
          put_Data_0_686 <= put_Data_0_659;
          put_size_680 <= 1;
          put_Data_1_690 <= put_Data_1_663;
          put_midKey_737 <= put_Key_1_660;
          put_Key_0_656 <= put_Key_2_664;
          put_Data_0_659 <= put_Data_2_667;
          put_Key_1_660 <= put_Key_3_668;
          put_Data_1_663 <= put_Data_3_671;
          put_size_653 <= 1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1166:<init>|  Btree.java:1165:splitLowButOne|  Btree.java:1756:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        423: begin
          put_root_738 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0076:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        424: begin
          put_freeNext_9_index_194 <= put_root_738;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1282:<init>|  Chip.java:1281:ExecuteTransaction|  Btree.java:0077:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        425: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0078:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        426: begin
          put_indexLeft_735 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0079:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        427: begin
          if (put_indexLeft_735 == 0) begin
            put_returnCode <= 20;
            put_stop <= 1;
          end
          put_isLeaf_740 <= 0;
          put_isFree_741 <= 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0082:<init>|  Btree.java:0081:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        428: begin
          put_freeNext_9_index_194 <= put_indexLeft_735;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          put_stuckIsLeaf_8_index_40 <= put_indexLeft_735;
          put_stuckIsLeaf_8_value_41 <= put_isLeaf_740;
          stuckIsLeaf_8_requestedAt <= step;
          stuckIsLeaf_8_finishedAt <= -1;
          put_stuckIsFree_11_index_197 <= put_indexLeft_735;
          put_stuckIsFree_11_value_198 <= put_isFree_741;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0097:<init>|  Btree.java:0096:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        429: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1289:<init>|  Chip.java:1288:waitResultOfTransaction|  Btree.java:0109:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        430: begin
          put_next_739 <= freeNext_freeNext_9_result_0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0110:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        431: begin
          put_freeNext_10_index_195 <= put_root_738;
          put_freeNext_10_value_196 <= put_next_739;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1345:<init>|  Chip.java:1344:ExecuteTransaction|  Btree.java:0111:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        432: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0112:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        433: begin
          if ((stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0113:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        434: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0114:allocate|  Btree.java:0152:allocateBranch|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        435: begin
          put_stuckSize_6_index_37 <= put_indexLeft_735;
          put_stuckSize_6_value_38 <= put_size_680;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_indexLeft_735;
          put_stuckKeys_2_value_26 <= put_Key_0_683;
          put_stuckKeys_2_value_27 <= put_Key_1_687;
          put_stuckKeys_2_value_28 <= put_Key_2_691;
          put_stuckKeys_2_value_29 <= put_Key_3_695;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_indexLeft_735;
          put_stuckData_4_value_32 <= put_Data_0_686;
          put_stuckData_4_value_33 <= put_Data_1_690;
          put_stuckData_4_value_34 <= put_Data_2_694;
          put_stuckData_4_value_35 <= put_Data_3_698;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        436: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        437: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        438: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1757:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        439: begin
          put_stuckSize_6_index_37 <= put_childData_734;
          put_stuckSize_6_value_38 <= put_size_653;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_childData_734;
          put_stuckKeys_2_value_26 <= put_Key_0_656;
          put_stuckKeys_2_value_27 <= put_Key_1_660;
          put_stuckKeys_2_value_28 <= put_Key_2_664;
          put_stuckKeys_2_value_29 <= put_Key_3_668;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_childData_734;
          put_stuckData_4_value_32 <= put_Data_0_659;
          put_stuckData_4_value_33 <= put_Data_1_663;
          put_stuckData_4_value_34 <= put_Data_2_667;
          put_stuckData_4_value_35 <= put_Data_3_671;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1758:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        440: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1758:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        441: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1758:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        442: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0336:stuckPut|  Btree.java:1758:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        443: begin
          case (put_size_626)
            0: begin
              put_Key_0_629 <= put_midKey_737;
              put_Data_0_632 <= put_indexLeft_735;
            end
            1: begin
              put_Key_1_633 <= put_midKey_737;
              put_Data_1_636 <= put_indexLeft_735;
            end
            2: begin
              put_Key_2_637 <= put_midKey_737;
              put_Data_2_640 <= put_indexLeft_735;
            end
            3: begin
              put_Key_3_641 <= put_midKey_737;
              put_Data_3_644 <= put_indexLeft_735;
            end
          endcase
          put_size_626 <= put_size_626+1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0424:<init>|  Btree.java:0423:Push|  Btree.java:1760:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        444: begin
          case (put_size_626)
            0: begin
              put_Key_0_629 <= put_midKey_737;
              put_Data_0_632 <= put_childData_734;
            end
            1: begin
              put_Key_1_633 <= put_midKey_737;
              put_Data_1_636 <= put_childData_734;
            end
            2: begin
              put_Key_2_637 <= put_midKey_737;
              put_Data_2_640 <= put_childData_734;
            end
            3: begin
              put_Key_3_641 <= put_midKey_737;
              put_Data_3_644 <= put_childData_734;
            end
          endcase
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0481:<init>|  Btree.java:0480:SetPastLastElement|  Btree.java:1761:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        445: begin
          put_stuckSize_6_index_37 <= put_index_625;
          put_stuckSize_6_value_38 <= put_size_626;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          put_stuckKeys_2_index_25 <= put_index_625;
          put_stuckKeys_2_value_26 <= put_Key_0_629;
          put_stuckKeys_2_value_27 <= put_Key_1_633;
          put_stuckKeys_2_value_28 <= put_Key_2_637;
          put_stuckKeys_2_value_29 <= put_Key_3_641;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          put_stuckData_4_index_31 <= put_index_625;
          put_stuckData_4_value_32 <= put_Data_0_632;
          put_stuckData_4_value_33 <= put_Data_1_636;
          put_stuckData_4_value_34 <= put_Data_2_640;
          put_stuckData_4_value_35 <= put_Data_3_644;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0314:<init>|  Btree.java:0313:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1762:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        446: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0328:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1762:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        447: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1762:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        448: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1352:<init>|  Chip.java:1351:waitResultOfTransaction|  Btree.java:0332:stuckPut|  Btree.java:0335:stuckPut|  Btree.java:1762:splitBranchAtTop|  Btree.java:2405:Else|  Chip.java:0620:<init>|  Btree.java:2401:<init>|  Btree.java:2400:Then|  Chip.java:0610:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        449: begin
          put_pc <= 451;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        450: begin
          put_parent_104 <= put_child_103;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2410:Else|  Chip.java:0620:<init>|  Btree.java:2399:<init>|  Btree.java:2398:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        451: begin
          put_pc <= 201;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:2414:Branch|  Btree.java:1414:code|  Chip.java:0530:<init>|  Btree.java:1389:<init>|  Btree.java:1388:<init>|  Btree.java:2376:<init>|  Btree.java:2375:code|  Chip.java:0530:<init>|  Btree.java:2360:<init>|  Btree.java:2359:code|  Chip.java:0530:<init>|  Btree.java:2334:<init>|  Btree.java:2333:put|  Btree.java:5942:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        452: begin
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:5945:<init>|  Btree.java:5944:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        453: begin
          put_l_3 <= put_k_0< 32 ? 1 : 0;
          put_pc <= put_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0788:<init>|  Chip.java:0788:Lt|  Btree.java:5950:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        454: begin
          if (put_l_3 >  0) begin
            put_pc <= 2;
          end
          else begin
            put_pc <= put_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0578:<init>|  Chip.java:0577:GONotZero|  Btree.java:5951:code|  Chip.java:0530:<init>|  Btree.java:5940:<init>|  Btree.java:5939:test_put_ascending|  Btree.java:7138:newTests|  Btree.java:7143:main|");
            $fclose(f);
          end
        end
        default: put_stop <= 1;
      endcase
    end
  end
  task chipPrint;
    begin
      integer o;
      o = $fopen("verilog/trace_verilog.txt", "a");
      if (!o) o = $fopen("../verilog/trace_verilog.txt", "a");
      if (!o) $display("Cannot create trace folder: verilog/trace_verilog.txt");
      $fwrite(o, "Chip: %-16s step: %1d, maxSteps: %1d, running: %1d\n", "Btree", step, maxSteps, !stop);
      $fwrite(o, "  Processes:\n");

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 0, "stuckIsLeaf", 1, stuckIsLeaf_pc, stuckIsLeaf_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsLeaf_memory[0]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[1]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[2]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[3]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[4]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[5]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[6]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[7]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[8]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[9]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[10]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[11]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[12]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[13]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[14]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[15]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[16]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[17]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[18]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[19]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[20]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[21]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[22]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[23]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[24]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[25]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[26]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[27]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[28]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[29]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[30]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckIsLeaf_7", stuckIsLeaf_7_requestedAt, stuckIsLeaf_7_finishedAt, stuckIsLeaf_stuckIsLeaf_7_returnCode, (stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step), (stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsLeaf_7_index_39", put_stuckIsLeaf_7_index_39);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsLeaf_8", stuckIsLeaf_8_requestedAt, stuckIsLeaf_8_finishedAt, stuckIsLeaf_stuckIsLeaf_8_returnCode, (stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step), (stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsLeaf_8_index_40", put_stuckIsLeaf_8_index_40);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsLeaf_8_value_41", put_stuckIsLeaf_8_value_41);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 1, "stuckIsFree", 1, stuckIsFree_pc, stuckIsFree_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsFree_memory[0]);
      $fwrite(o, ", %2d", stuckIsFree_memory[1]);
      $fwrite(o, ", %2d", stuckIsFree_memory[2]);
      $fwrite(o, ", %2d", stuckIsFree_memory[3]);
      $fwrite(o, ", %2d", stuckIsFree_memory[4]);
      $fwrite(o, ", %2d", stuckIsFree_memory[5]);
      $fwrite(o, ", %2d", stuckIsFree_memory[6]);
      $fwrite(o, ", %2d", stuckIsFree_memory[7]);
      $fwrite(o, ", %2d", stuckIsFree_memory[8]);
      $fwrite(o, ", %2d", stuckIsFree_memory[9]);
      $fwrite(o, ", %2d", stuckIsFree_memory[10]);
      $fwrite(o, ", %2d", stuckIsFree_memory[11]);
      $fwrite(o, ", %2d", stuckIsFree_memory[12]);
      $fwrite(o, ", %2d", stuckIsFree_memory[13]);
      $fwrite(o, ", %2d", stuckIsFree_memory[14]);
      $fwrite(o, ", %2d", stuckIsFree_memory[15]);
      $fwrite(o, ", %2d", stuckIsFree_memory[16]);
      $fwrite(o, ", %2d", stuckIsFree_memory[17]);
      $fwrite(o, ", %2d", stuckIsFree_memory[18]);
      $fwrite(o, ", %2d", stuckIsFree_memory[19]);
      $fwrite(o, ", %2d", stuckIsFree_memory[20]);
      $fwrite(o, ", %2d", stuckIsFree_memory[21]);
      $fwrite(o, ", %2d", stuckIsFree_memory[22]);
      $fwrite(o, ", %2d", stuckIsFree_memory[23]);
      $fwrite(o, ", %2d", stuckIsFree_memory[24]);
      $fwrite(o, ", %2d", stuckIsFree_memory[25]);
      $fwrite(o, ", %2d", stuckIsFree_memory[26]);
      $fwrite(o, ", %2d", stuckIsFree_memory[27]);
      $fwrite(o, ", %2d", stuckIsFree_memory[28]);
      $fwrite(o, ", %2d", stuckIsFree_memory[29]);
      $fwrite(o, ", %2d", stuckIsFree_memory[30]);
      $fwrite(o, ", %2d", stuckIsFree_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsFree_11", stuckIsFree_11_requestedAt, stuckIsFree_11_finishedAt, stuckIsFree_stuckIsFree_11_returnCode, (stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step), (stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsFree_11_index_197", put_stuckIsFree_11_index_197);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckIsFree_11_value_198", put_stuckIsFree_11_value_198);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 2, "freeNext", 1, freeNext_pc, freeNext_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 6, 1);
      $fwrite(o, "        %2d", freeNext_memory[0]);
      $fwrite(o, ", %2d", freeNext_memory[1]);
      $fwrite(o, ", %2d", freeNext_memory[2]);
      $fwrite(o, ", %2d", freeNext_memory[3]);
      $fwrite(o, ", %2d", freeNext_memory[4]);
      $fwrite(o, ", %2d", freeNext_memory[5]);
      $fwrite(o, ", %2d", freeNext_memory[6]);
      $fwrite(o, ", %2d", freeNext_memory[7]);
      $fwrite(o, ", %2d", freeNext_memory[8]);
      $fwrite(o, ", %2d", freeNext_memory[9]);
      $fwrite(o, ", %2d", freeNext_memory[10]);
      $fwrite(o, ", %2d", freeNext_memory[11]);
      $fwrite(o, ", %2d", freeNext_memory[12]);
      $fwrite(o, ", %2d", freeNext_memory[13]);
      $fwrite(o, ", %2d", freeNext_memory[14]);
      $fwrite(o, ", %2d", freeNext_memory[15]);
      $fwrite(o, ", %2d", freeNext_memory[16]);
      $fwrite(o, ", %2d", freeNext_memory[17]);
      $fwrite(o, ", %2d", freeNext_memory[18]);
      $fwrite(o, ", %2d", freeNext_memory[19]);
      $fwrite(o, ", %2d", freeNext_memory[20]);
      $fwrite(o, ", %2d", freeNext_memory[21]);
      $fwrite(o, ", %2d", freeNext_memory[22]);
      $fwrite(o, ", %2d", freeNext_memory[23]);
      $fwrite(o, ", %2d", freeNext_memory[24]);
      $fwrite(o, ", %2d", freeNext_memory[25]);
      $fwrite(o, ", %2d", freeNext_memory[26]);
      $fwrite(o, ", %2d", freeNext_memory[27]);
      $fwrite(o, ", %2d", freeNext_memory[28]);
      $fwrite(o, ", %2d", freeNext_memory[29]);
      $fwrite(o, ", %2d", freeNext_memory[30]);
      $fwrite(o, ", %2d", freeNext_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "freeNext_9", freeNext_9_requestedAt, freeNext_9_finishedAt, freeNext_freeNext_9_returnCode, (freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step), (freeNext_9_requestedAt < freeNext_9_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_freeNext_9_index_194", put_freeNext_9_index_194);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "freeNext_10", freeNext_10_requestedAt, freeNext_10_finishedAt, freeNext_freeNext_10_returnCode, (freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step), (freeNext_10_requestedAt < freeNext_10_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_freeNext_10_index_195", put_freeNext_10_index_195);

      $fwrite(o, "            %-38s = %1d\n", "put_freeNext_10_value_196", put_freeNext_10_value_196);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 3, "stuckSize", 1, stuckSize_pc, stuckSize_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 3, 1);
      $fwrite(o, "        %2d", stuckSize_memory[0]);
      $fwrite(o, ", %2d", stuckSize_memory[1]);
      $fwrite(o, ", %2d", stuckSize_memory[2]);
      $fwrite(o, ", %2d", stuckSize_memory[3]);
      $fwrite(o, ", %2d", stuckSize_memory[4]);
      $fwrite(o, ", %2d", stuckSize_memory[5]);
      $fwrite(o, ", %2d", stuckSize_memory[6]);
      $fwrite(o, ", %2d", stuckSize_memory[7]);
      $fwrite(o, ", %2d", stuckSize_memory[8]);
      $fwrite(o, ", %2d", stuckSize_memory[9]);
      $fwrite(o, ", %2d", stuckSize_memory[10]);
      $fwrite(o, ", %2d", stuckSize_memory[11]);
      $fwrite(o, ", %2d", stuckSize_memory[12]);
      $fwrite(o, ", %2d", stuckSize_memory[13]);
      $fwrite(o, ", %2d", stuckSize_memory[14]);
      $fwrite(o, ", %2d", stuckSize_memory[15]);
      $fwrite(o, ", %2d", stuckSize_memory[16]);
      $fwrite(o, ", %2d", stuckSize_memory[17]);
      $fwrite(o, ", %2d", stuckSize_memory[18]);
      $fwrite(o, ", %2d", stuckSize_memory[19]);
      $fwrite(o, ", %2d", stuckSize_memory[20]);
      $fwrite(o, ", %2d", stuckSize_memory[21]);
      $fwrite(o, ", %2d", stuckSize_memory[22]);
      $fwrite(o, ", %2d", stuckSize_memory[23]);
      $fwrite(o, ", %2d", stuckSize_memory[24]);
      $fwrite(o, ", %2d", stuckSize_memory[25]);
      $fwrite(o, ", %2d", stuckSize_memory[26]);
      $fwrite(o, ", %2d", stuckSize_memory[27]);
      $fwrite(o, ", %2d", stuckSize_memory[28]);
      $fwrite(o, ", %2d", stuckSize_memory[29]);
      $fwrite(o, ", %2d", stuckSize_memory[30]);
      $fwrite(o, ", %2d", stuckSize_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckSize_5", stuckSize_5_requestedAt, stuckSize_5_finishedAt, stuckSize_stuckSize_5_returnCode, (stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step), (stuckSize_5_requestedAt < stuckSize_5_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckSize_5_index_36", put_stuckSize_5_index_36);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckSize_6", stuckSize_6_requestedAt, stuckSize_6_finishedAt, stuckSize_stuckSize_6_returnCode, (stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step), (stuckSize_6_requestedAt < stuckSize_6_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckSize_6_index_37", put_stuckSize_6_index_37);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckSize_6_value_38", put_stuckSize_6_value_38);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 4, "stuckKeys", 1, stuckKeys_pc, stuckKeys_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckKeys_memory[0]);
      $fwrite(o, ", %2d", stuckKeys_memory[1]);
      $fwrite(o, ", %2d", stuckKeys_memory[2]);
      $fwrite(o, ", %2d", stuckKeys_memory[3]);
      $fwrite(o, ", %2d", stuckKeys_memory[4]);
      $fwrite(o, ", %2d", stuckKeys_memory[5]);
      $fwrite(o, ", %2d", stuckKeys_memory[6]);
      $fwrite(o, ", %2d", stuckKeys_memory[7]);
      $fwrite(o, ", %2d", stuckKeys_memory[8]);
      $fwrite(o, ", %2d", stuckKeys_memory[9]);
      $fwrite(o, ", %2d", stuckKeys_memory[10]);
      $fwrite(o, ", %2d", stuckKeys_memory[11]);
      $fwrite(o, ", %2d", stuckKeys_memory[12]);
      $fwrite(o, ", %2d", stuckKeys_memory[13]);
      $fwrite(o, ", %2d", stuckKeys_memory[14]);
      $fwrite(o, ", %2d", stuckKeys_memory[15]);
      $fwrite(o, ", %2d", stuckKeys_memory[16]);
      $fwrite(o, ", %2d", stuckKeys_memory[17]);
      $fwrite(o, ", %2d", stuckKeys_memory[18]);
      $fwrite(o, ", %2d", stuckKeys_memory[19]);
      $fwrite(o, ", %2d", stuckKeys_memory[20]);
      $fwrite(o, ", %2d", stuckKeys_memory[21]);
      $fwrite(o, ", %2d", stuckKeys_memory[22]);
      $fwrite(o, ", %2d", stuckKeys_memory[23]);
      $fwrite(o, ", %2d", stuckKeys_memory[24]);
      $fwrite(o, ", %2d", stuckKeys_memory[25]);
      $fwrite(o, ", %2d", stuckKeys_memory[26]);
      $fwrite(o, ", %2d", stuckKeys_memory[27]);
      $fwrite(o, ", %2d", stuckKeys_memory[28]);
      $fwrite(o, ", %2d", stuckKeys_memory[29]);
      $fwrite(o, ", %2d", stuckKeys_memory[30]);
      $fwrite(o, ", %2d", stuckKeys_memory[31]);
      $fwrite(o, ", %2d", stuckKeys_memory[32]);
      $fwrite(o, ", %2d", stuckKeys_memory[33]);
      $fwrite(o, ", %2d", stuckKeys_memory[34]);
      $fwrite(o, ", %2d", stuckKeys_memory[35]);
      $fwrite(o, ", %2d", stuckKeys_memory[36]);
      $fwrite(o, ", %2d", stuckKeys_memory[37]);
      $fwrite(o, ", %2d", stuckKeys_memory[38]);
      $fwrite(o, ", %2d", stuckKeys_memory[39]);
      $fwrite(o, ", %2d", stuckKeys_memory[40]);
      $fwrite(o, ", %2d", stuckKeys_memory[41]);
      $fwrite(o, ", %2d", stuckKeys_memory[42]);
      $fwrite(o, ", %2d", stuckKeys_memory[43]);
      $fwrite(o, ", %2d", stuckKeys_memory[44]);
      $fwrite(o, ", %2d", stuckKeys_memory[45]);
      $fwrite(o, ", %2d", stuckKeys_memory[46]);
      $fwrite(o, ", %2d", stuckKeys_memory[47]);
      $fwrite(o, ", %2d", stuckKeys_memory[48]);
      $fwrite(o, ", %2d", stuckKeys_memory[49]);
      $fwrite(o, ", %2d", stuckKeys_memory[50]);
      $fwrite(o, ", %2d", stuckKeys_memory[51]);
      $fwrite(o, ", %2d", stuckKeys_memory[52]);
      $fwrite(o, ", %2d", stuckKeys_memory[53]);
      $fwrite(o, ", %2d", stuckKeys_memory[54]);
      $fwrite(o, ", %2d", stuckKeys_memory[55]);
      $fwrite(o, ", %2d", stuckKeys_memory[56]);
      $fwrite(o, ", %2d", stuckKeys_memory[57]);
      $fwrite(o, ", %2d", stuckKeys_memory[58]);
      $fwrite(o, ", %2d", stuckKeys_memory[59]);
      $fwrite(o, ", %2d", stuckKeys_memory[60]);
      $fwrite(o, ", %2d", stuckKeys_memory[61]);
      $fwrite(o, ", %2d", stuckKeys_memory[62]);
      $fwrite(o, ", %2d", stuckKeys_memory[63]);
      $fwrite(o, ", %2d", stuckKeys_memory[64]);
      $fwrite(o, ", %2d", stuckKeys_memory[65]);
      $fwrite(o, ", %2d", stuckKeys_memory[66]);
      $fwrite(o, ", %2d", stuckKeys_memory[67]);
      $fwrite(o, ", %2d", stuckKeys_memory[68]);
      $fwrite(o, ", %2d", stuckKeys_memory[69]);
      $fwrite(o, ", %2d", stuckKeys_memory[70]);
      $fwrite(o, ", %2d", stuckKeys_memory[71]);
      $fwrite(o, ", %2d", stuckKeys_memory[72]);
      $fwrite(o, ", %2d", stuckKeys_memory[73]);
      $fwrite(o, ", %2d", stuckKeys_memory[74]);
      $fwrite(o, ", %2d", stuckKeys_memory[75]);
      $fwrite(o, ", %2d", stuckKeys_memory[76]);
      $fwrite(o, ", %2d", stuckKeys_memory[77]);
      $fwrite(o, ", %2d", stuckKeys_memory[78]);
      $fwrite(o, ", %2d", stuckKeys_memory[79]);
      $fwrite(o, ", %2d", stuckKeys_memory[80]);
      $fwrite(o, ", %2d", stuckKeys_memory[81]);
      $fwrite(o, ", %2d", stuckKeys_memory[82]);
      $fwrite(o, ", %2d", stuckKeys_memory[83]);
      $fwrite(o, ", %2d", stuckKeys_memory[84]);
      $fwrite(o, ", %2d", stuckKeys_memory[85]);
      $fwrite(o, ", %2d", stuckKeys_memory[86]);
      $fwrite(o, ", %2d", stuckKeys_memory[87]);
      $fwrite(o, ", %2d", stuckKeys_memory[88]);
      $fwrite(o, ", %2d", stuckKeys_memory[89]);
      $fwrite(o, ", %2d", stuckKeys_memory[90]);
      $fwrite(o, ", %2d", stuckKeys_memory[91]);
      $fwrite(o, ", %2d", stuckKeys_memory[92]);
      $fwrite(o, ", %2d", stuckKeys_memory[93]);
      $fwrite(o, ", %2d", stuckKeys_memory[94]);
      $fwrite(o, ", %2d", stuckKeys_memory[95]);
      $fwrite(o, ", %2d", stuckKeys_memory[96]);
      $fwrite(o, ", %2d", stuckKeys_memory[97]);
      $fwrite(o, ", %2d", stuckKeys_memory[98]);
      $fwrite(o, ", %2d", stuckKeys_memory[99]);
      $fwrite(o, ", %2d", stuckKeys_memory[100]);
      $fwrite(o, ", %2d", stuckKeys_memory[101]);
      $fwrite(o, ", %2d", stuckKeys_memory[102]);
      $fwrite(o, ", %2d", stuckKeys_memory[103]);
      $fwrite(o, ", %2d", stuckKeys_memory[104]);
      $fwrite(o, ", %2d", stuckKeys_memory[105]);
      $fwrite(o, ", %2d", stuckKeys_memory[106]);
      $fwrite(o, ", %2d", stuckKeys_memory[107]);
      $fwrite(o, ", %2d", stuckKeys_memory[108]);
      $fwrite(o, ", %2d", stuckKeys_memory[109]);
      $fwrite(o, ", %2d", stuckKeys_memory[110]);
      $fwrite(o, ", %2d", stuckKeys_memory[111]);
      $fwrite(o, ", %2d", stuckKeys_memory[112]);
      $fwrite(o, ", %2d", stuckKeys_memory[113]);
      $fwrite(o, ", %2d", stuckKeys_memory[114]);
      $fwrite(o, ", %2d", stuckKeys_memory[115]);
      $fwrite(o, ", %2d", stuckKeys_memory[116]);
      $fwrite(o, ", %2d", stuckKeys_memory[117]);
      $fwrite(o, ", %2d", stuckKeys_memory[118]);
      $fwrite(o, ", %2d", stuckKeys_memory[119]);
      $fwrite(o, ", %2d", stuckKeys_memory[120]);
      $fwrite(o, ", %2d", stuckKeys_memory[121]);
      $fwrite(o, ", %2d", stuckKeys_memory[122]);
      $fwrite(o, ", %2d", stuckKeys_memory[123]);
      $fwrite(o, ", %2d", stuckKeys_memory[124]);
      $fwrite(o, ", %2d", stuckKeys_memory[125]);
      $fwrite(o, ", %2d", stuckKeys_memory[126]);
      $fwrite(o, ", %2d", stuckKeys_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckKeys_1", stuckKeys_1_requestedAt, stuckKeys_1_finishedAt, stuckKeys_stuckKeys_1_returnCode, (stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step), (stuckKeys_1_requestedAt < stuckKeys_1_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_1_index_24", put_stuckKeys_1_index_24);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckKeys_2", stuckKeys_2_requestedAt, stuckKeys_2_finishedAt, stuckKeys_stuckKeys_2_returnCode, (stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step), (stuckKeys_2_requestedAt < stuckKeys_2_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_index_25", put_stuckKeys_2_index_25);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_26", put_stuckKeys_2_value_26);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_27", put_stuckKeys_2_value_27);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_28", put_stuckKeys_2_value_28);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckKeys_2_value_29", put_stuckKeys_2_value_29);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 5, "stuckData", 1, stuckData_pc, stuckData_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckData_memory[0]);
      $fwrite(o, ", %2d", stuckData_memory[1]);
      $fwrite(o, ", %2d", stuckData_memory[2]);
      $fwrite(o, ", %2d", stuckData_memory[3]);
      $fwrite(o, ", %2d", stuckData_memory[4]);
      $fwrite(o, ", %2d", stuckData_memory[5]);
      $fwrite(o, ", %2d", stuckData_memory[6]);
      $fwrite(o, ", %2d", stuckData_memory[7]);
      $fwrite(o, ", %2d", stuckData_memory[8]);
      $fwrite(o, ", %2d", stuckData_memory[9]);
      $fwrite(o, ", %2d", stuckData_memory[10]);
      $fwrite(o, ", %2d", stuckData_memory[11]);
      $fwrite(o, ", %2d", stuckData_memory[12]);
      $fwrite(o, ", %2d", stuckData_memory[13]);
      $fwrite(o, ", %2d", stuckData_memory[14]);
      $fwrite(o, ", %2d", stuckData_memory[15]);
      $fwrite(o, ", %2d", stuckData_memory[16]);
      $fwrite(o, ", %2d", stuckData_memory[17]);
      $fwrite(o, ", %2d", stuckData_memory[18]);
      $fwrite(o, ", %2d", stuckData_memory[19]);
      $fwrite(o, ", %2d", stuckData_memory[20]);
      $fwrite(o, ", %2d", stuckData_memory[21]);
      $fwrite(o, ", %2d", stuckData_memory[22]);
      $fwrite(o, ", %2d", stuckData_memory[23]);
      $fwrite(o, ", %2d", stuckData_memory[24]);
      $fwrite(o, ", %2d", stuckData_memory[25]);
      $fwrite(o, ", %2d", stuckData_memory[26]);
      $fwrite(o, ", %2d", stuckData_memory[27]);
      $fwrite(o, ", %2d", stuckData_memory[28]);
      $fwrite(o, ", %2d", stuckData_memory[29]);
      $fwrite(o, ", %2d", stuckData_memory[30]);
      $fwrite(o, ", %2d", stuckData_memory[31]);
      $fwrite(o, ", %2d", stuckData_memory[32]);
      $fwrite(o, ", %2d", stuckData_memory[33]);
      $fwrite(o, ", %2d", stuckData_memory[34]);
      $fwrite(o, ", %2d", stuckData_memory[35]);
      $fwrite(o, ", %2d", stuckData_memory[36]);
      $fwrite(o, ", %2d", stuckData_memory[37]);
      $fwrite(o, ", %2d", stuckData_memory[38]);
      $fwrite(o, ", %2d", stuckData_memory[39]);
      $fwrite(o, ", %2d", stuckData_memory[40]);
      $fwrite(o, ", %2d", stuckData_memory[41]);
      $fwrite(o, ", %2d", stuckData_memory[42]);
      $fwrite(o, ", %2d", stuckData_memory[43]);
      $fwrite(o, ", %2d", stuckData_memory[44]);
      $fwrite(o, ", %2d", stuckData_memory[45]);
      $fwrite(o, ", %2d", stuckData_memory[46]);
      $fwrite(o, ", %2d", stuckData_memory[47]);
      $fwrite(o, ", %2d", stuckData_memory[48]);
      $fwrite(o, ", %2d", stuckData_memory[49]);
      $fwrite(o, ", %2d", stuckData_memory[50]);
      $fwrite(o, ", %2d", stuckData_memory[51]);
      $fwrite(o, ", %2d", stuckData_memory[52]);
      $fwrite(o, ", %2d", stuckData_memory[53]);
      $fwrite(o, ", %2d", stuckData_memory[54]);
      $fwrite(o, ", %2d", stuckData_memory[55]);
      $fwrite(o, ", %2d", stuckData_memory[56]);
      $fwrite(o, ", %2d", stuckData_memory[57]);
      $fwrite(o, ", %2d", stuckData_memory[58]);
      $fwrite(o, ", %2d", stuckData_memory[59]);
      $fwrite(o, ", %2d", stuckData_memory[60]);
      $fwrite(o, ", %2d", stuckData_memory[61]);
      $fwrite(o, ", %2d", stuckData_memory[62]);
      $fwrite(o, ", %2d", stuckData_memory[63]);
      $fwrite(o, ", %2d", stuckData_memory[64]);
      $fwrite(o, ", %2d", stuckData_memory[65]);
      $fwrite(o, ", %2d", stuckData_memory[66]);
      $fwrite(o, ", %2d", stuckData_memory[67]);
      $fwrite(o, ", %2d", stuckData_memory[68]);
      $fwrite(o, ", %2d", stuckData_memory[69]);
      $fwrite(o, ", %2d", stuckData_memory[70]);
      $fwrite(o, ", %2d", stuckData_memory[71]);
      $fwrite(o, ", %2d", stuckData_memory[72]);
      $fwrite(o, ", %2d", stuckData_memory[73]);
      $fwrite(o, ", %2d", stuckData_memory[74]);
      $fwrite(o, ", %2d", stuckData_memory[75]);
      $fwrite(o, ", %2d", stuckData_memory[76]);
      $fwrite(o, ", %2d", stuckData_memory[77]);
      $fwrite(o, ", %2d", stuckData_memory[78]);
      $fwrite(o, ", %2d", stuckData_memory[79]);
      $fwrite(o, ", %2d", stuckData_memory[80]);
      $fwrite(o, ", %2d", stuckData_memory[81]);
      $fwrite(o, ", %2d", stuckData_memory[82]);
      $fwrite(o, ", %2d", stuckData_memory[83]);
      $fwrite(o, ", %2d", stuckData_memory[84]);
      $fwrite(o, ", %2d", stuckData_memory[85]);
      $fwrite(o, ", %2d", stuckData_memory[86]);
      $fwrite(o, ", %2d", stuckData_memory[87]);
      $fwrite(o, ", %2d", stuckData_memory[88]);
      $fwrite(o, ", %2d", stuckData_memory[89]);
      $fwrite(o, ", %2d", stuckData_memory[90]);
      $fwrite(o, ", %2d", stuckData_memory[91]);
      $fwrite(o, ", %2d", stuckData_memory[92]);
      $fwrite(o, ", %2d", stuckData_memory[93]);
      $fwrite(o, ", %2d", stuckData_memory[94]);
      $fwrite(o, ", %2d", stuckData_memory[95]);
      $fwrite(o, ", %2d", stuckData_memory[96]);
      $fwrite(o, ", %2d", stuckData_memory[97]);
      $fwrite(o, ", %2d", stuckData_memory[98]);
      $fwrite(o, ", %2d", stuckData_memory[99]);
      $fwrite(o, ", %2d", stuckData_memory[100]);
      $fwrite(o, ", %2d", stuckData_memory[101]);
      $fwrite(o, ", %2d", stuckData_memory[102]);
      $fwrite(o, ", %2d", stuckData_memory[103]);
      $fwrite(o, ", %2d", stuckData_memory[104]);
      $fwrite(o, ", %2d", stuckData_memory[105]);
      $fwrite(o, ", %2d", stuckData_memory[106]);
      $fwrite(o, ", %2d", stuckData_memory[107]);
      $fwrite(o, ", %2d", stuckData_memory[108]);
      $fwrite(o, ", %2d", stuckData_memory[109]);
      $fwrite(o, ", %2d", stuckData_memory[110]);
      $fwrite(o, ", %2d", stuckData_memory[111]);
      $fwrite(o, ", %2d", stuckData_memory[112]);
      $fwrite(o, ", %2d", stuckData_memory[113]);
      $fwrite(o, ", %2d", stuckData_memory[114]);
      $fwrite(o, ", %2d", stuckData_memory[115]);
      $fwrite(o, ", %2d", stuckData_memory[116]);
      $fwrite(o, ", %2d", stuckData_memory[117]);
      $fwrite(o, ", %2d", stuckData_memory[118]);
      $fwrite(o, ", %2d", stuckData_memory[119]);
      $fwrite(o, ", %2d", stuckData_memory[120]);
      $fwrite(o, ", %2d", stuckData_memory[121]);
      $fwrite(o, ", %2d", stuckData_memory[122]);
      $fwrite(o, ", %2d", stuckData_memory[123]);
      $fwrite(o, ", %2d", stuckData_memory[124]);
      $fwrite(o, ", %2d", stuckData_memory[125]);
      $fwrite(o, ", %2d", stuckData_memory[126]);
      $fwrite(o, ", %2d", stuckData_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckData_3", stuckData_3_requestedAt, stuckData_3_finishedAt, stuckData_stuckData_3_returnCode, (stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step), (stuckData_3_requestedAt < stuckData_3_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_3_index_30", put_stuckData_3_index_30);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckData_4", stuckData_4_requestedAt, stuckData_4_finishedAt, stuckData_stuckData_4_returnCode, (stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step), (stuckData_4_requestedAt < stuckData_4_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_index_31", put_stuckData_4_index_31);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_32", put_stuckData_4_value_32);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_33", put_stuckData_4_value_33);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_34", put_stuckData_4_value_34);

      $fwrite(o, "            %-38s = %1d\n", "put_stuckData_4_value_35", put_stuckData_4_value_35);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 6, "put", 455, put_pc, put_returnCode);
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_k_0", put_k_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_d_1", put_d_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_2", put_i_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_l_3", put_l_3);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_4", put_index_4);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_5", put_size_5);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_6", put_isLeaf_6);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_7", put_nextFree_7);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_8", put_Key_0_8);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_9", put_KeyCompares_0_9);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_10", put_KeyCollapse_0_10);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_11", put_Data_0_11);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_12", put_Key_1_12);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_13", put_KeyCompares_1_13);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_14", put_KeyCollapse_1_14);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_15", put_Data_1_15);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_16", put_Key_2_16);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_17", put_KeyCompares_2_17);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_18", put_KeyCollapse_2_18);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_19", put_Data_2_19);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_20", put_Key_3_20);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_21", put_KeyCompares_3_21);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_22", put_KeyCollapse_3_22);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_23", put_Data_3_23);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_1_index_24", put_stuckKeys_1_index_24);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_index_25", put_stuckKeys_2_index_25);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_26", put_stuckKeys_2_value_26);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_27", put_stuckKeys_2_value_27);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_28", put_stuckKeys_2_value_28);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckKeys_2_value_29", put_stuckKeys_2_value_29);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_3_index_30", put_stuckData_3_index_30);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_index_31", put_stuckData_4_index_31);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_32", put_stuckData_4_value_32);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_33", put_stuckData_4_value_33);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_34", put_stuckData_4_value_34);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckData_4_value_35", put_stuckData_4_value_35);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckSize_5_index_36", put_stuckSize_5_index_36);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckSize_6_index_37", put_stuckSize_6_index_37);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckSize_6_value_38", put_stuckSize_6_value_38);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsLeaf_7_index_39", put_stuckIsLeaf_7_index_39);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsLeaf_8_index_40", put_stuckIsLeaf_8_index_40);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsLeaf_8_value_41", put_stuckIsLeaf_8_value_41);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_42", put_Found_42);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_43", put_Key_43);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_44", put_FoundKey_44);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_45", put_Data_45);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_46", put_BtreeIndex_46);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_47", put_StuckIndex_47);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_48", put_MergeSuccess_48);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_49", put_index_49);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_50", put_size_50);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_51", put_isLeaf_51);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_52", put_nextFree_52);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_53", put_Key_0_53);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_54", put_KeyCompares_0_54);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_55", put_KeyCollapse_0_55);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_56", put_Data_0_56);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_57", put_Key_1_57);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_58", put_KeyCompares_1_58);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_59", put_KeyCollapse_1_59);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_60", put_Data_1_60);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_61", put_Key_2_61);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_62", put_KeyCompares_2_62);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_63", put_KeyCollapse_2_63);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_64", put_Data_2_64);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_65", put_Key_3_65);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_66", put_KeyCompares_3_66);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_67", put_KeyCollapse_3_67);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_68", put_Data_3_68);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_69", put_Found_69);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_70", put_Key_70);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_71", put_FoundKey_71);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_72", put_Data_72);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_73", put_BtreeIndex_73);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_74", put_StuckIndex_74);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_75", put_MergeSuccess_75);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_76", put_index_76);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_77", put_size_77);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_78", put_isLeaf_78);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_79", put_nextFree_79);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_80", put_Key_0_80);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_81", put_KeyCompares_0_81);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_82", put_KeyCollapse_0_82);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_83", put_Data_0_83);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_84", put_Key_1_84);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_85", put_KeyCompares_1_85);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_86", put_KeyCollapse_1_86);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_87", put_Data_1_87);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_88", put_Key_2_88);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_89", put_KeyCompares_2_89);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_90", put_KeyCollapse_2_90);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_91", put_Data_2_91);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_92", put_Key_3_92);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_93", put_KeyCompares_3_93);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_94", put_KeyCollapse_3_94);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_95", put_Data_3_95);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_96", put_Found_96);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_97", put_Key_97);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_98", put_FoundKey_98);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_99", put_Data_99);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_100", put_BtreeIndex_100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_101", put_StuckIndex_101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_102", put_MergeSuccess_102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_child_103", put_child_103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_parent_104", put_parent_104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childInparent_105", put_childInparent_105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_found_106", put_found_106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_full_107", put_full_107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_108", put_i_108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_notFull_109", put_notFull_109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_110", put_index_110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_111", put_size_111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_112", put_isLeaf_112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_113", put_nextFree_113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_114", put_Key_0_114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_115", put_KeyCompares_0_115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_116", put_KeyCollapse_0_116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_117", put_Data_0_117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_118", put_Key_1_118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_119", put_KeyCompares_1_119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_120", put_KeyCollapse_1_120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_121", put_Data_1_121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_122", put_Key_2_122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_123", put_KeyCompares_2_123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_124", put_KeyCollapse_2_124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_125", put_Data_2_125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_126", put_Key_3_126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_127", put_KeyCompares_3_127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_128", put_KeyCollapse_3_128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_129", put_Data_3_129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_130", put_Found_130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_131", put_Key_131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_132", put_FoundKey_132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_133", put_Data_133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_134", put_BtreeIndex_134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_135", put_StuckIndex_135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_136", put_MergeSuccess_136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_137", put_index_137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_138", put_size_138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_139", put_isLeaf_139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_140", put_nextFree_140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_141", put_Key_0_141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_142", put_KeyCompares_0_142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_143", put_KeyCollapse_0_143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_144", put_Data_0_144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_145", put_Key_1_145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_146", put_KeyCompares_1_146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_147", put_KeyCollapse_1_147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_148", put_Data_1_148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_149", put_Key_2_149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_150", put_KeyCompares_2_150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_151", put_KeyCollapse_2_151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_152", put_Data_2_152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_153", put_Key_3_153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_154", put_KeyCompares_3_154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_155", put_KeyCollapse_3_155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_156", put_Data_3_156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_157", put_Found_157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_158", put_Key_158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_159", put_FoundKey_159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_160", put_Data_160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_161", put_BtreeIndex_161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_162", put_StuckIndex_162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_163", put_MergeSuccess_163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_164", put_index_164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_165", put_size_165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_166", put_isLeaf_166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_167", put_nextFree_167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_168", put_Key_0_168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_169", put_KeyCompares_0_169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_170", put_KeyCollapse_0_170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_171", put_Data_0_171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_172", put_Key_1_172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_173", put_KeyCompares_1_173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_174", put_KeyCollapse_1_174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_175", put_Data_1_175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_176", put_Key_2_176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_177", put_KeyCompares_2_177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_178", put_KeyCollapse_2_178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_179", put_Data_2_179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_180", put_Key_3_180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_181", put_KeyCompares_3_181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_182", put_KeyCollapse_3_182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_183", put_Data_3_183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_184", put_Found_184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_185", put_Key_185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_186", put_FoundKey_186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_187", put_Data_187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_188", put_BtreeIndex_188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_189", put_StuckIndex_189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_190", put_MergeSuccess_190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_191", put_indexLeft_191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_192", put_indexRight_192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_193", put_midKey_193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_freeNext_9_index_194", put_freeNext_9_index_194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_freeNext_10_index_195", put_freeNext_10_index_195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_freeNext_10_value_196", put_freeNext_10_value_196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsFree_11_index_197", put_stuckIsFree_11_index_197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_stuckIsFree_11_value_198", put_stuckIsFree_11_value_198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_199", put_root_199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_200", put_next_200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_201", put_isLeaf_201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_202", put_isFree_202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_203", put_root_203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_204", put_next_204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_205", put_isLeaf_205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_206", put_isFree_206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_207", put_i_207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_notFull_208", put_notFull_208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_209", put_index_209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_210", put_size_210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_211", put_isLeaf_211);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_212", put_nextFree_212);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_213", put_Key_0_213);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_214", put_KeyCompares_0_214);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_215", put_KeyCollapse_0_215);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_216", put_Data_0_216);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_217", put_Key_1_217);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_218", put_KeyCompares_1_218);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_219", put_KeyCollapse_1_219);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_220", put_Data_1_220);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_221", put_Key_2_221);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_222", put_KeyCompares_2_222);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_223", put_KeyCollapse_2_223);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_224", put_Data_2_224);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_225", put_Key_3_225);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_226", put_KeyCompares_3_226);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_227", put_KeyCollapse_3_227);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_228", put_Data_3_228);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_229", put_Found_229);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_230", put_Key_230);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_231", put_FoundKey_231);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_232", put_Data_232);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_233", put_BtreeIndex_233);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_234", put_StuckIndex_234);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_235", put_MergeSuccess_235);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_236", put_index_236);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_237", put_size_237);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_238", put_isLeaf_238);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_239", put_nextFree_239);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_240", put_Key_0_240);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_241", put_KeyCompares_0_241);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_242", put_KeyCollapse_0_242);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_243", put_Data_0_243);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_244", put_Key_1_244);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_245", put_KeyCompares_1_245);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_246", put_KeyCollapse_1_246);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_247", put_Data_1_247);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_248", put_Key_2_248);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_249", put_KeyCompares_2_249);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_250", put_KeyCollapse_2_250);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_251", put_Data_2_251);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_252", put_Key_3_252);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_253", put_KeyCompares_3_253);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_254", put_KeyCollapse_3_254);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_255", put_Data_3_255);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_256", put_Found_256);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_257", put_Key_257);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_258", put_FoundKey_258);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_259", put_Data_259);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_260", put_BtreeIndex_260);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_261", put_StuckIndex_261);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_262", put_MergeSuccess_262);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_263", put_index_263);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_264", put_size_264);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_265", put_isLeaf_265);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_266", put_nextFree_266);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_267", put_Key_0_267);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_268", put_KeyCompares_0_268);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_269", put_KeyCollapse_0_269);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_270", put_Data_0_270);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_271", put_Key_1_271);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_272", put_KeyCompares_1_272);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_273", put_KeyCollapse_1_273);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_274", put_Data_1_274);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_275", put_Key_2_275);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_276", put_KeyCompares_2_276);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_277", put_KeyCollapse_2_277);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_278", put_Data_2_278);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_279", put_Key_3_279);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_280", put_KeyCompares_3_280);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_281", put_KeyCollapse_3_281);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_282", put_Data_3_282);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_283", put_Found_283);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_284", put_Key_284);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_285", put_FoundKey_285);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_286", put_Data_286);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_287", put_BtreeIndex_287);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_288", put_StuckIndex_288);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_289", put_MergeSuccess_289);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_290", put_indexLeft_290);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_291", put_indexRight_291);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_292", put_midKey_292);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_293", put_root_293);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_294", put_next_294);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_295", put_isLeaf_295);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_296", put_isFree_296);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_297", put_root_297);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_298", put_next_298);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_299", put_isLeaf_299);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_300", put_isFree_300);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_301", put_index_301);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_302", put_size_302);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_303", put_isLeaf_303);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_304", put_nextFree_304);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_305", put_Key_0_305);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_306", put_KeyCompares_0_306);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_307", put_KeyCollapse_0_307);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_308", put_Data_0_308);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_309", put_Key_1_309);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_310", put_KeyCompares_1_310);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_311", put_KeyCollapse_1_311);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_312", put_Data_1_312);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_313", put_Key_2_313);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_314", put_KeyCompares_2_314);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_315", put_KeyCollapse_2_315);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_316", put_Data_2_316);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_317", put_Key_3_317);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_318", put_KeyCompares_3_318);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_319", put_KeyCollapse_3_319);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_320", put_Data_3_320);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_321", put_Found_321);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_322", put_Key_322);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_323", put_FoundKey_323);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_324", put_Data_324);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_325", put_BtreeIndex_325);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_326", put_StuckIndex_326);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_327", put_MergeSuccess_327);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_328", put_index_328);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_329", put_size_329);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_330", put_isLeaf_330);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_331", put_nextFree_331);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_332", put_Key_0_332);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_333", put_KeyCompares_0_333);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_334", put_KeyCollapse_0_334);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_335", put_Data_0_335);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_336", put_Key_1_336);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_337", put_KeyCompares_1_337);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_338", put_KeyCollapse_1_338);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_339", put_Data_1_339);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_340", put_Key_2_340);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_341", put_KeyCompares_2_341);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_342", put_KeyCollapse_2_342);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_343", put_Data_2_343);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_344", put_Key_3_344);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_345", put_KeyCompares_3_345);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_346", put_KeyCollapse_3_346);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_347", put_Data_3_347);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_348", put_Found_348);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_349", put_Key_349);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_350", put_FoundKey_350);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_351", put_Data_351);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_352", put_BtreeIndex_352);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_353", put_StuckIndex_353);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_354", put_MergeSuccess_354);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_355", put_index_355);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_356", put_size_356);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_357", put_isLeaf_357);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_358", put_nextFree_358);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_359", put_Key_0_359);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_360", put_KeyCompares_0_360);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_361", put_KeyCollapse_0_361);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_362", put_Data_0_362);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_363", put_Key_1_363);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_364", put_KeyCompares_1_364);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_365", put_KeyCollapse_1_365);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_366", put_Data_1_366);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_367", put_Key_2_367);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_368", put_KeyCompares_2_368);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_369", put_KeyCollapse_2_369);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_370", put_Data_2_370);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_371", put_Key_3_371);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_372", put_KeyCompares_3_372);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_373", put_KeyCollapse_3_373);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_374", put_Data_3_374);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_375", put_Found_375);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_376", put_Key_376);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_377", put_FoundKey_377);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_378", put_Data_378);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_379", put_BtreeIndex_379);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_380", put_StuckIndex_380);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_381", put_MergeSuccess_381);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_382", put_index_382);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_383", put_size_383);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_384", put_isLeaf_384);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_385", put_nextFree_385);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_386", put_Key_0_386);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_387", put_KeyCompares_0_387);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_388", put_KeyCollapse_0_388);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_389", put_Data_0_389);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_390", put_Key_1_390);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_391", put_KeyCompares_1_391);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_392", put_KeyCollapse_1_392);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_393", put_Data_1_393);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_394", put_Key_2_394);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_395", put_KeyCompares_2_395);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_396", put_KeyCollapse_2_396);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_397", put_Data_2_397);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_398", put_Key_3_398);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_399", put_KeyCompares_3_399);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_400", put_KeyCollapse_3_400);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_401", put_Data_3_401);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_402", put_Found_402);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_403", put_Key_403);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_404", put_FoundKey_404);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_405", put_Data_405);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_406", put_BtreeIndex_406);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_407", put_StuckIndex_407);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_408", put_MergeSuccess_408);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_409", put_childKey_409);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_410", put_childData_410);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_411", put_indexLeft_411);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_412", put_indexRight_412);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_413", put_midKey_413);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_414", put_root_414);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_415", put_next_415);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_416", put_isLeaf_416);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_417", put_isFree_417);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_418", put_index_418);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_419", put_size_419);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_420", put_isLeaf_420);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_421", put_nextFree_421);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_422", put_Key_0_422);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_423", put_KeyCompares_0_423);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_424", put_KeyCollapse_0_424);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_425", put_Data_0_425);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_426", put_Key_1_426);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_427", put_KeyCompares_1_427);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_428", put_KeyCollapse_1_428);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_429", put_Data_1_429);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_430", put_Key_2_430);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_431", put_KeyCompares_2_431);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_432", put_KeyCollapse_2_432);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_433", put_Data_2_433);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_434", put_Key_3_434);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_435", put_KeyCompares_3_435);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_436", put_KeyCollapse_3_436);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_437", put_Data_3_437);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_438", put_Found_438);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_439", put_Key_439);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_440", put_FoundKey_440);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_441", put_Data_441);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_442", put_BtreeIndex_442);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_443", put_StuckIndex_443);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_444", put_MergeSuccess_444);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_445", put_index_445);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_446", put_size_446);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_447", put_isLeaf_447);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_448", put_nextFree_448);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_449", put_Key_0_449);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_450", put_KeyCompares_0_450);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_451", put_KeyCollapse_0_451);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_452", put_Data_0_452);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_453", put_Key_1_453);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_454", put_KeyCompares_1_454);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_455", put_KeyCollapse_1_455);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_456", put_Data_1_456);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_457", put_Key_2_457);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_458", put_KeyCompares_2_458);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_459", put_KeyCollapse_2_459);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_460", put_Data_2_460);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_461", put_Key_3_461);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_462", put_KeyCompares_3_462);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_463", put_KeyCollapse_3_463);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_464", put_Data_3_464);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_465", put_Found_465);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_466", put_Key_466);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_467", put_FoundKey_467);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_468", put_Data_468);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_469", put_BtreeIndex_469);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_470", put_StuckIndex_470);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_471", put_MergeSuccess_471);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_472", put_index_472);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_473", put_size_473);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_474", put_isLeaf_474);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_475", put_nextFree_475);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_476", put_Key_0_476);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_477", put_KeyCompares_0_477);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_478", put_KeyCollapse_0_478);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_479", put_Data_0_479);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_480", put_Key_1_480);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_481", put_KeyCompares_1_481);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_482", put_KeyCollapse_1_482);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_483", put_Data_1_483);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_484", put_Key_2_484);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_485", put_KeyCompares_2_485);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_486", put_KeyCollapse_2_486);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_487", put_Data_2_487);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_488", put_Key_3_488);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_489", put_KeyCompares_3_489);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_490", put_KeyCollapse_3_490);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_491", put_Data_3_491);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_492", put_Found_492);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_493", put_Key_493);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_494", put_FoundKey_494);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_495", put_Data_495);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_496", put_BtreeIndex_496);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_497", put_StuckIndex_497);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_498", put_MergeSuccess_498);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childIndex_499", put_childIndex_499);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_leftIndex_500", put_leftIndex_500);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_501", put_midKey_501);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_502", put_root_502);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_503", put_next_503);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_504", put_isLeaf_504);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_505", put_isFree_505);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_i_506", put_i_506);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_notFull_507", put_notFull_507);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_508", put_index_508);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_509", put_size_509);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_510", put_isLeaf_510);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_511", put_nextFree_511);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_512", put_Key_0_512);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_513", put_KeyCompares_0_513);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_514", put_KeyCollapse_0_514);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_515", put_Data_0_515);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_516", put_Key_1_516);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_517", put_KeyCompares_1_517);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_518", put_KeyCollapse_1_518);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_519", put_Data_1_519);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_520", put_Key_2_520);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_521", put_KeyCompares_2_521);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_522", put_KeyCollapse_2_522);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_523", put_Data_2_523);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_524", put_Key_3_524);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_525", put_KeyCompares_3_525);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_526", put_KeyCollapse_3_526);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_527", put_Data_3_527);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_528", put_Found_528);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_529", put_Key_529);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_530", put_FoundKey_530);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_531", put_Data_531);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_532", put_BtreeIndex_532);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_533", put_StuckIndex_533);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_534", put_MergeSuccess_534);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_535", put_index_535);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_536", put_size_536);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_537", put_isLeaf_537);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_538", put_nextFree_538);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_539", put_Key_0_539);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_540", put_KeyCompares_0_540);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_541", put_KeyCollapse_0_541);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_542", put_Data_0_542);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_543", put_Key_1_543);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_544", put_KeyCompares_1_544);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_545", put_KeyCollapse_1_545);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_546", put_Data_1_546);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_547", put_Key_2_547);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_548", put_KeyCompares_2_548);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_549", put_KeyCollapse_2_549);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_550", put_Data_2_550);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_551", put_Key_3_551);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_552", put_KeyCompares_3_552);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_553", put_KeyCollapse_3_553);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_554", put_Data_3_554);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_555", put_Found_555);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_556", put_Key_556);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_557", put_FoundKey_557);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_558", put_Data_558);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_559", put_BtreeIndex_559);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_560", put_StuckIndex_560);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_561", put_MergeSuccess_561);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_562", put_index_562);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_563", put_size_563);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_564", put_isLeaf_564);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_565", put_nextFree_565);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_566", put_Key_0_566);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_567", put_KeyCompares_0_567);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_568", put_KeyCollapse_0_568);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_569", put_Data_0_569);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_570", put_Key_1_570);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_571", put_KeyCompares_1_571);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_572", put_KeyCollapse_1_572);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_573", put_Data_1_573);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_574", put_Key_2_574);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_575", put_KeyCompares_2_575);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_576", put_KeyCollapse_2_576);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_577", put_Data_2_577);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_578", put_Key_3_578);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_579", put_KeyCompares_3_579);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_580", put_KeyCollapse_3_580);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_581", put_Data_3_581);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_582", put_Found_582);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_583", put_Key_583);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_584", put_FoundKey_584);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_585", put_Data_585);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_586", put_BtreeIndex_586);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_587", put_StuckIndex_587);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_588", put_MergeSuccess_588);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_589", put_index_589);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_590", put_size_590);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_591", put_isLeaf_591);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_592", put_nextFree_592);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_593", put_Key_0_593);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_594", put_KeyCompares_0_594);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_595", put_KeyCollapse_0_595);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_596", put_Data_0_596);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_597", put_Key_1_597);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_598", put_KeyCompares_1_598);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_599", put_KeyCollapse_1_599);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_600", put_Data_1_600);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_601", put_Key_2_601);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_602", put_KeyCompares_2_602);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_603", put_KeyCollapse_2_603);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_604", put_Data_2_604);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_605", put_Key_3_605);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_606", put_KeyCompares_3_606);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_607", put_KeyCollapse_3_607);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_608", put_Data_3_608);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_609", put_Found_609);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_610", put_Key_610);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_611", put_FoundKey_611);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_612", put_Data_612);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_613", put_BtreeIndex_613);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_614", put_StuckIndex_614);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_615", put_MergeSuccess_615);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_616", put_childKey_616);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_617", put_childData_617);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_618", put_indexLeft_618);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_619", put_indexRight_619);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_620", put_midKey_620);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_621", put_root_621);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_622", put_next_622);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_623", put_isLeaf_623);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_624", put_isFree_624);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_625", put_index_625);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_626", put_size_626);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_627", put_isLeaf_627);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_628", put_nextFree_628);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_629", put_Key_0_629);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_630", put_KeyCompares_0_630);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_631", put_KeyCollapse_0_631);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_632", put_Data_0_632);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_633", put_Key_1_633);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_634", put_KeyCompares_1_634);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_635", put_KeyCollapse_1_635);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_636", put_Data_1_636);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_637", put_Key_2_637);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_638", put_KeyCompares_2_638);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_639", put_KeyCollapse_2_639);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_640", put_Data_2_640);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_641", put_Key_3_641);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_642", put_KeyCompares_3_642);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_643", put_KeyCollapse_3_643);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_644", put_Data_3_644);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_645", put_Found_645);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_646", put_Key_646);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_647", put_FoundKey_647);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_648", put_Data_648);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_649", put_BtreeIndex_649);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_650", put_StuckIndex_650);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_651", put_MergeSuccess_651);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_652", put_index_652);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_653", put_size_653);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_654", put_isLeaf_654);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_655", put_nextFree_655);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_656", put_Key_0_656);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_657", put_KeyCompares_0_657);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_658", put_KeyCollapse_0_658);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_659", put_Data_0_659);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_660", put_Key_1_660);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_661", put_KeyCompares_1_661);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_662", put_KeyCollapse_1_662);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_663", put_Data_1_663);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_664", put_Key_2_664);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_665", put_KeyCompares_2_665);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_666", put_KeyCollapse_2_666);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_667", put_Data_2_667);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_668", put_Key_3_668);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_669", put_KeyCompares_3_669);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_670", put_KeyCollapse_3_670);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_671", put_Data_3_671);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_672", put_Found_672);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_673", put_Key_673);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_674", put_FoundKey_674);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_675", put_Data_675);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_676", put_BtreeIndex_676);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_677", put_StuckIndex_677);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_678", put_MergeSuccess_678);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_679", put_index_679);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_680", put_size_680);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_681", put_isLeaf_681);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_682", put_nextFree_682);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_683", put_Key_0_683);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_684", put_KeyCompares_0_684);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_685", put_KeyCollapse_0_685);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_686", put_Data_0_686);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_687", put_Key_1_687);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_688", put_KeyCompares_1_688);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_689", put_KeyCollapse_1_689);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_690", put_Data_1_690);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_691", put_Key_2_691);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_692", put_KeyCompares_2_692);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_693", put_KeyCollapse_2_693);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_694", put_Data_2_694);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_695", put_Key_3_695);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_696", put_KeyCompares_3_696);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_697", put_KeyCollapse_3_697);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_698", put_Data_3_698);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_699", put_Found_699);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_700", put_Key_700);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_701", put_FoundKey_701);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_702", put_Data_702);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_703", put_BtreeIndex_703);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_704", put_StuckIndex_704);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_705", put_MergeSuccess_705);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_index_706", put_index_706);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_size_707", put_size_707);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_708", put_isLeaf_708);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_nextFree_709", put_nextFree_709);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_0_710", put_Key_0_710);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_0_711", put_KeyCompares_0_711);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_0_712", put_KeyCollapse_0_712);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_0_713", put_Data_0_713);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_1_714", put_Key_1_714);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_1_715", put_KeyCompares_1_715);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_1_716", put_KeyCollapse_1_716);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_1_717", put_Data_1_717);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_2_718", put_Key_2_718);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_2_719", put_KeyCompares_2_719);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_2_720", put_KeyCollapse_2_720);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_2_721", put_Data_2_721);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_3_722", put_Key_3_722);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCompares_3_723", put_KeyCompares_3_723);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_KeyCollapse_3_724", put_KeyCollapse_3_724);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_3_725", put_Data_3_725);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Found_726", put_Found_726);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Key_727", put_Key_727);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_FoundKey_728", put_FoundKey_728);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_Data_729", put_Data_729);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_BtreeIndex_730", put_BtreeIndex_730);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_StuckIndex_731", put_StuckIndex_731);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_MergeSuccess_732", put_MergeSuccess_732);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childKey_733", put_childKey_733);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_childData_734", put_childData_734);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexLeft_735", put_indexLeft_735);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_indexRight_736", put_indexRight_736);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_midKey_737", put_midKey_737);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_root_738", put_root_738);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_next_739", put_next_739);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isLeaf_740", put_isLeaf_740);
      $fwrite(o, "        Register: %-32s = %1d\n",  "put_isFree_741", put_isFree_741);
      $fclose(o);
    end
  endtask
endmodule
