//-----------------------------------------------------------------------------
// Database on a chip test bench
// Philip R Brenan at appaapps dot com, Appa Apps Ltd Inc., 2025
//------------------------------------------------------------------------------
`timescale 10ps/1ps
module Btree;                                                                      // Test bench for database on a chip
  reg                    stop;                                                  // Program has stopped when this goes high
  reg                   clock;                                                  // Clock
  integer                step;                                                  // Step of the simulation
  integer            maxSteps;                                                  // Maximum number of steps to execute
  integer          returnCode;                                                  // Return code
  integer      processCurrent;                                                  // To ensure we get the same results in Java and Verilog we have to run the processes single threaded in a constant order

  assign stop = stuckIsLeaf_stop||stuckIsFree_stop||freeNext_stop||stuckSize_stop||stuckKeys_stop||stuckData_stop||findAndInsert_stop;                                                             // Or of process stop fields

  initial begin
    returnCode = 0;
    maxSteps = 2000;
    for(step = -1; step < 0 || step < maxSteps && !stop; step = step + 1) begin // Steps below zero are run unconditionally to initialize each process so that Java and Verilog start in sync at step zero

      processCurrent = 0; clock = 0; #1; clock = 1; #1; // process_stuckIsLeaf_0000
      processCurrent = 1; clock = 0; #1; clock = 1; #1; // process_stuckIsFree_0001
      processCurrent = 2; clock = 0; #1; clock = 1; #1; // process_freeNext_0002
      processCurrent = 3; clock = 0; #1; clock = 1; #1; // process_stuckSize_0003
      processCurrent = 4; clock = 0; #1; clock = 1; #1; // process_stuckKeys_0004
      processCurrent = 5; clock = 0; #1; clock = 1; #1; // process_stuckData_0005
      processCurrent = 6; clock = 0; #1; clock = 1; #1; // process_findAndInsert_0006
      if (step >= 0) chipPrint();                                            // Steps prior to zero are for initialization to make Java and Verilog match
    end
    if (!stop) $finish(1); else $finish(0);                                // Set return code depending on whether the simulation halted
  end
  // Process: stuckIsLeaf  process_stuckIsLeaf_0000
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsLeaf_memory[32*1];
  reg [1-1:0] stuckIsLeaf_stuckIsLeaf_7_result_0;
  integer stuckIsLeaf_7_requestedAt;
  integer stuckIsLeaf_7_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_7_returnCode;
  integer stuckIsLeaf_8_requestedAt;
  integer stuckIsLeaf_8_finishedAt;
  integer stuckIsLeaf_stuckIsLeaf_8_returnCode;
  integer stuckIsLeaf_pc;
  integer stuckIsLeaf_stop;
  integer stuckIsLeaf_returnCode;
  integer stuckIsLeaf_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsLeaf_pc <= 0;
      stuckIsLeaf_stop <= 0;
      stuckIsLeaf_returnCode <= 0;
      stuckIsLeaf_stuckIsLeaf_7_result_0 <= 0;
      stuckIsLeaf_7_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_7_returnCode <= 0;
      stuckIsLeaf_8_finishedAt <= -1;
      stuckIsLeaf_stuckIsLeaf_8_returnCode <= 0;
      for(stuckIsLeaf_memory_index = 0; stuckIsLeaf_memory_index < 1; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
      stuckIsLeaf_memory[1] <= 1;
      stuckIsLeaf_memory[2] <= 1;
      stuckIsLeaf_memory[3] <= 1;
      stuckIsLeaf_memory[4] <= 1;
      for(stuckIsLeaf_memory_index = 5; stuckIsLeaf_memory_index < 7; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
      stuckIsLeaf_memory[7] <= 1;
      stuckIsLeaf_memory[8] <= 1;
      stuckIsLeaf_memory[9] <= 1;
      stuckIsLeaf_memory[10] <= 1;
      for(stuckIsLeaf_memory_index = 11; stuckIsLeaf_memory_index < 12; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
      stuckIsLeaf_memory[12] <= 1;
      for(stuckIsLeaf_memory_index = 13; stuckIsLeaf_memory_index < 32; stuckIsLeaf_memory_index = stuckIsLeaf_memory_index + 1) stuckIsLeaf_memory[stuckIsLeaf_memory_index] <= 0;
    end
    else if (processCurrent == 0) begin
      case(stuckIsLeaf_pc)
        0: begin
          if ((stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step)) begin
            stuckIsLeaf_stuckIsLeaf_7_result_0 <= stuckIsLeaf_memory[findAndInsert_stuckIsLeaf_7_index_35*1+0];
            stuckIsLeaf_7_finishedAt <= step;
          end
          else if ((stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step)) begin
            stuckIsLeaf_memory[findAndInsert_stuckIsLeaf_8_index_36*1+0] <= findAndInsert_stuckIsLeaf_8_value_37;
            stuckIsLeaf_8_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsLeaf_stop <= 1;
      endcase
    end
  end
  // Process: stuckIsFree  process_stuckIsFree_0001
  (* ram_style = "block" *)
  reg [1-1:0] stuckIsFree_memory[32*1];
  integer stuckIsFree_11_requestedAt;
  integer stuckIsFree_11_finishedAt;
  integer stuckIsFree_stuckIsFree_11_returnCode;
  integer stuckIsFree_pc;
  integer stuckIsFree_stop;
  integer stuckIsFree_returnCode;
  integer stuckIsFree_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckIsFree_pc <= 0;
      stuckIsFree_stop <= 0;
      stuckIsFree_returnCode <= 0;
      stuckIsFree_11_finishedAt <= -1;
      stuckIsFree_stuckIsFree_11_returnCode <= 0;
      for(stuckIsFree_memory_index = 0; stuckIsFree_memory_index < 12; stuckIsFree_memory_index = stuckIsFree_memory_index + 1) stuckIsFree_memory[stuckIsFree_memory_index] <= 0;
      stuckIsFree_memory[12] <= 1;
      stuckIsFree_memory[13] <= 1;
      stuckIsFree_memory[14] <= 1;
      stuckIsFree_memory[15] <= 1;
      stuckIsFree_memory[16] <= 1;
      stuckIsFree_memory[17] <= 1;
      stuckIsFree_memory[18] <= 1;
      stuckIsFree_memory[19] <= 1;
      stuckIsFree_memory[20] <= 1;
      stuckIsFree_memory[21] <= 1;
      stuckIsFree_memory[22] <= 1;
      stuckIsFree_memory[23] <= 1;
      stuckIsFree_memory[24] <= 1;
      stuckIsFree_memory[25] <= 1;
      stuckIsFree_memory[26] <= 1;
      stuckIsFree_memory[27] <= 1;
      stuckIsFree_memory[28] <= 1;
      stuckIsFree_memory[29] <= 1;
      stuckIsFree_memory[30] <= 1;
      stuckIsFree_memory[31] <= 1;
    end
    else if (processCurrent == 1) begin
      case(stuckIsFree_pc)
        0: begin
          if ((stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step)) begin
            stuckIsFree_memory[findAndInsert_stuckIsFree_11_index_163*1+0] <= findAndInsert_stuckIsFree_11_value_164;
            stuckIsFree_11_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckIsFree_stop <= 1;
      endcase
    end
  end
  // Process: freeNext  process_freeNext_0002
  (* ram_style = "block" *)
  reg [6-1:0] freeNext_memory[32*1];
  reg [6-1:0] freeNext_freeNext_9_result_0;
  integer freeNext_9_requestedAt;
  integer freeNext_9_finishedAt;
  integer freeNext_freeNext_9_returnCode;
  integer freeNext_10_requestedAt;
  integer freeNext_10_finishedAt;
  integer freeNext_freeNext_10_returnCode;
  integer freeNext_pc;
  integer freeNext_stop;
  integer freeNext_returnCode;
  integer freeNext_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      freeNext_pc <= 0;
      freeNext_stop <= 0;
      freeNext_returnCode <= 0;
      freeNext_freeNext_9_result_0 <= 0;
      freeNext_9_finishedAt <= -1;
      freeNext_freeNext_9_returnCode <= 0;
      freeNext_10_finishedAt <= -1;
      freeNext_freeNext_10_returnCode <= 0;
      freeNext_memory[0] <= 12;
      freeNext_memory[1] <= 2;
      freeNext_memory[2] <= 3;
      freeNext_memory[3] <= 4;
      freeNext_memory[4] <= 5;
      freeNext_memory[5] <= 6;
      freeNext_memory[6] <= 12;
      freeNext_memory[7] <= 8;
      freeNext_memory[8] <= 9;
      freeNext_memory[9] <= 11;
      freeNext_memory[10] <= 9;
      freeNext_memory[11] <= 12;
      freeNext_memory[12] <= 13;
      freeNext_memory[13] <= 14;
      freeNext_memory[14] <= 15;
      freeNext_memory[15] <= 16;
      freeNext_memory[16] <= 17;
      freeNext_memory[17] <= 18;
      freeNext_memory[18] <= 19;
      freeNext_memory[19] <= 20;
      freeNext_memory[20] <= 21;
      freeNext_memory[21] <= 22;
      freeNext_memory[22] <= 23;
      freeNext_memory[23] <= 24;
      freeNext_memory[24] <= 25;
      freeNext_memory[25] <= 26;
      freeNext_memory[26] <= 27;
      freeNext_memory[27] <= 28;
      freeNext_memory[28] <= 29;
      freeNext_memory[29] <= 30;
      freeNext_memory[30] <= 31;
      for(freeNext_memory_index = 31; freeNext_memory_index < 32; freeNext_memory_index = freeNext_memory_index + 1) freeNext_memory[freeNext_memory_index] <= 0;
    end
    else if (processCurrent == 2) begin
      case(freeNext_pc)
        0: begin
          if ((freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step)) begin
            freeNext_freeNext_9_result_0 <= freeNext_memory[findAndInsert_freeNext_9_index_160*1+0];
            freeNext_9_finishedAt <= step;
          end
          else if ((freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step)) begin
            freeNext_memory[findAndInsert_freeNext_10_index_161*1+0] <= findAndInsert_freeNext_10_value_162;
            freeNext_10_finishedAt <= step;
          end
          else begin
          end
        end
        default: freeNext_stop <= 1;
      endcase
    end
  end
  // Process: stuckSize  process_stuckSize_0003
  (* ram_style = "block" *)
  reg [3-1:0] stuckSize_memory[32*1];
  reg [3-1:0] stuckSize_stuckSize_5_result_0;
  integer stuckSize_5_requestedAt;
  integer stuckSize_5_finishedAt;
  integer stuckSize_stuckSize_5_returnCode;
  integer stuckSize_6_requestedAt;
  integer stuckSize_6_finishedAt;
  integer stuckSize_stuckSize_6_returnCode;
  integer stuckSize_pc;
  integer stuckSize_stop;
  integer stuckSize_returnCode;
  integer stuckSize_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckSize_pc <= 0;
      stuckSize_stop <= 0;
      stuckSize_returnCode <= 0;
      stuckSize_stuckSize_5_result_0 <= 0;
      stuckSize_5_finishedAt <= -1;
      stuckSize_stuckSize_5_returnCode <= 0;
      stuckSize_6_finishedAt <= -1;
      stuckSize_stuckSize_6_returnCode <= 0;
      stuckSize_memory[0] <= 2;
      stuckSize_memory[1] <= 4;
      stuckSize_memory[2] <= 4;
      stuckSize_memory[3] <= 4;
      stuckSize_memory[4] <= 4;
      stuckSize_memory[5] <= 3;
      stuckSize_memory[6] <= 1;
      stuckSize_memory[7] <= 4;
      stuckSize_memory[8] <= 4;
      stuckSize_memory[9] <= 4;
      stuckSize_memory[10] <= 4;
      stuckSize_memory[11] <= 1;
      stuckSize_memory[12] <= 2;
      for(stuckSize_memory_index = 13; stuckSize_memory_index < 32; stuckSize_memory_index = stuckSize_memory_index + 1) stuckSize_memory[stuckSize_memory_index] <= 0;
    end
    else if (processCurrent == 3) begin
      case(stuckSize_pc)
        0: begin
          if ((stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step)) begin
            stuckSize_stuckSize_5_result_0 <= stuckSize_memory[findAndInsert_stuckSize_5_index_32*1+0];
            stuckSize_5_finishedAt <= step;
          end
          else if ((stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step)) begin
            stuckSize_memory[findAndInsert_stuckSize_6_index_33*1+0] <= findAndInsert_stuckSize_6_value_34;
            stuckSize_6_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckSize_stop <= 1;
      endcase
    end
  end
  // Process: stuckKeys  process_stuckKeys_0004
  (* ram_style = "block" *)
  reg [8-1:0] stuckKeys_memory[32*4];
  reg [8-1:0] stuckKeys_stuckKeys_1_result_0;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_1;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_2;
  reg [8-1:0] stuckKeys_stuckKeys_1_result_3;
  integer stuckKeys_1_requestedAt;
  integer stuckKeys_1_finishedAt;
  integer stuckKeys_stuckKeys_1_returnCode;
  integer stuckKeys_2_requestedAt;
  integer stuckKeys_2_finishedAt;
  integer stuckKeys_stuckKeys_2_returnCode;
  integer stuckKeys_pc;
  integer stuckKeys_stop;
  integer stuckKeys_returnCode;
  integer stuckKeys_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckKeys_pc <= 0;
      stuckKeys_stop <= 0;
      stuckKeys_returnCode <= 0;
      stuckKeys_stuckKeys_1_result_0 <= 0;
      stuckKeys_stuckKeys_1_result_1 <= 0;
      stuckKeys_stuckKeys_1_result_2 <= 0;
      stuckKeys_stuckKeys_1_result_3 <= 0;
      stuckKeys_1_finishedAt <= -1;
      stuckKeys_stuckKeys_1_returnCode <= 0;
      stuckKeys_2_finishedAt <= -1;
      stuckKeys_stuckKeys_2_returnCode <= 0;
      stuckKeys_memory[0] <= 16;
      stuckKeys_memory[1] <= 24;
      stuckKeys_memory[2] <= 24;
      stuckKeys_memory[3] <= 10;
      stuckKeys_memory[4] <= 1;
      stuckKeys_memory[5] <= 2;
      stuckKeys_memory[6] <= 3;
      stuckKeys_memory[7] <= 4;
      stuckKeys_memory[8] <= 29;
      stuckKeys_memory[9] <= 30;
      stuckKeys_memory[10] <= 31;
      stuckKeys_memory[11] <= 32;
      stuckKeys_memory[12] <= 5;
      stuckKeys_memory[13] <= 6;
      stuckKeys_memory[14] <= 7;
      stuckKeys_memory[15] <= 8;
      stuckKeys_memory[16] <= 9;
      stuckKeys_memory[17] <= 10;
      stuckKeys_memory[18] <= 11;
      stuckKeys_memory[19] <= 12;
      stuckKeys_memory[20] <= 4;
      stuckKeys_memory[21] <= 8;
      stuckKeys_memory[22] <= 12;
      for(stuckKeys_memory_index = 23; stuckKeys_memory_index < 24; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
      stuckKeys_memory[24] <= 20;
      for(stuckKeys_memory_index = 25; stuckKeys_memory_index < 28; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
      stuckKeys_memory[28] <= 13;
      stuckKeys_memory[29] <= 14;
      stuckKeys_memory[30] <= 15;
      stuckKeys_memory[31] <= 16;
      stuckKeys_memory[32] <= 17;
      stuckKeys_memory[33] <= 18;
      stuckKeys_memory[34] <= 19;
      stuckKeys_memory[35] <= 20;
      stuckKeys_memory[36] <= 25;
      stuckKeys_memory[37] <= 26;
      stuckKeys_memory[38] <= 27;
      stuckKeys_memory[39] <= 28;
      stuckKeys_memory[40] <= 21;
      stuckKeys_memory[41] <= 22;
      stuckKeys_memory[42] <= 23;
      stuckKeys_memory[43] <= 24;
      stuckKeys_memory[44] <= 28;
      for(stuckKeys_memory_index = 45; stuckKeys_memory_index < 46; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
      stuckKeys_memory[46] <= 28;
      for(stuckKeys_memory_index = 47; stuckKeys_memory_index < 48; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
      stuckKeys_memory[48] <= 27;
      stuckKeys_memory[49] <= 28;
      for(stuckKeys_memory_index = 50; stuckKeys_memory_index < 128; stuckKeys_memory_index = stuckKeys_memory_index + 1) stuckKeys_memory[stuckKeys_memory_index] <= 0;
    end
    else if (processCurrent == 4) begin
      case(stuckKeys_pc)
        0: begin
          if ((stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step)) begin
            stuckKeys_stuckKeys_1_result_0 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+0];
            stuckKeys_stuckKeys_1_result_1 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+1];
            stuckKeys_stuckKeys_1_result_2 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+2];
            stuckKeys_stuckKeys_1_result_3 <= stuckKeys_memory[findAndInsert_stuckKeys_1_index_20*4+3];
            stuckKeys_1_finishedAt <= step;
          end
          else if ((stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step)) begin
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+0] <= findAndInsert_stuckKeys_2_value_22;
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+1] <= findAndInsert_stuckKeys_2_value_23;
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+2] <= findAndInsert_stuckKeys_2_value_24;
            stuckKeys_memory[findAndInsert_stuckKeys_2_index_21*4+3] <= findAndInsert_stuckKeys_2_value_25;
            stuckKeys_2_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckKeys_stop <= 1;
      endcase
    end
  end
  // Process: stuckData  process_stuckData_0005
  (* ram_style = "block" *)
  reg [8-1:0] stuckData_memory[32*4];
  reg [8-1:0] stuckData_stuckData_3_result_0;
  reg [8-1:0] stuckData_stuckData_3_result_1;
  reg [8-1:0] stuckData_stuckData_3_result_2;
  reg [8-1:0] stuckData_stuckData_3_result_3;
  integer stuckData_3_requestedAt;
  integer stuckData_3_finishedAt;
  integer stuckData_stuckData_3_returnCode;
  integer stuckData_4_requestedAt;
  integer stuckData_4_finishedAt;
  integer stuckData_stuckData_4_returnCode;
  integer stuckData_pc;
  integer stuckData_stop;
  integer stuckData_returnCode;
  integer stuckData_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      stuckData_pc <= 0;
      stuckData_stop <= 0;
      stuckData_returnCode <= 0;
      stuckData_stuckData_3_result_0 <= 0;
      stuckData_stuckData_3_result_1 <= 0;
      stuckData_stuckData_3_result_2 <= 0;
      stuckData_stuckData_3_result_3 <= 0;
      stuckData_3_finishedAt <= -1;
      stuckData_stuckData_3_returnCode <= 0;
      stuckData_4_finishedAt <= -1;
      stuckData_stuckData_4_returnCode <= 0;
      stuckData_memory[0] <= 5;
      stuckData_memory[1] <= 6;
      stuckData_memory[2] <= 11;
      stuckData_memory[3] <= 2;
      stuckData_memory[4] <= 2;
      stuckData_memory[5] <= 3;
      stuckData_memory[6] <= 4;
      stuckData_memory[7] <= 5;
      stuckData_memory[8] <= 30;
      stuckData_memory[9] <= 31;
      stuckData_memory[10] <= 32;
      stuckData_memory[11] <= 33;
      stuckData_memory[12] <= 6;
      stuckData_memory[13] <= 7;
      stuckData_memory[14] <= 8;
      stuckData_memory[15] <= 9;
      stuckData_memory[16] <= 10;
      stuckData_memory[17] <= 11;
      stuckData_memory[18] <= 12;
      stuckData_memory[19] <= 13;
      stuckData_memory[20] <= 1;
      stuckData_memory[21] <= 3;
      stuckData_memory[22] <= 4;
      stuckData_memory[23] <= 7;
      stuckData_memory[24] <= 8;
      stuckData_memory[25] <= 10;
      for(stuckData_memory_index = 26; stuckData_memory_index < 28; stuckData_memory_index = stuckData_memory_index + 1) stuckData_memory[stuckData_memory_index] <= 0;
      stuckData_memory[28] <= 14;
      stuckData_memory[29] <= 15;
      stuckData_memory[30] <= 16;
      stuckData_memory[31] <= 17;
      stuckData_memory[32] <= 18;
      stuckData_memory[33] <= 19;
      stuckData_memory[34] <= 20;
      stuckData_memory[35] <= 21;
      stuckData_memory[36] <= 26;
      stuckData_memory[37] <= 27;
      stuckData_memory[38] <= 28;
      stuckData_memory[39] <= 29;
      stuckData_memory[40] <= 22;
      stuckData_memory[41] <= 23;
      stuckData_memory[42] <= 24;
      stuckData_memory[43] <= 25;
      stuckData_memory[44] <= 9;
      stuckData_memory[45] <= 2;
      stuckData_memory[46] <= 9;
      stuckData_memory[47] <= 2;
      stuckData_memory[48] <= 28;
      stuckData_memory[49] <= 29;
      for(stuckData_memory_index = 50; stuckData_memory_index < 128; stuckData_memory_index = stuckData_memory_index + 1) stuckData_memory[stuckData_memory_index] <= 0;
    end
    else if (processCurrent == 5) begin
      case(stuckData_pc)
        0: begin
          if ((stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step)) begin
            stuckData_stuckData_3_result_0 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+0];
            stuckData_stuckData_3_result_1 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+1];
            stuckData_stuckData_3_result_2 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+2];
            stuckData_stuckData_3_result_3 <= stuckData_memory[findAndInsert_stuckData_3_index_26*4+3];
            stuckData_3_finishedAt <= step;
          end
          else if ((stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step)) begin
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+0] <= findAndInsert_stuckData_4_value_28;
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+1] <= findAndInsert_stuckData_4_value_29;
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+2] <= findAndInsert_stuckData_4_value_30;
            stuckData_memory[findAndInsert_stuckData_4_index_27*4+3] <= findAndInsert_stuckData_4_value_31;
            stuckData_4_finishedAt <= step;
          end
          else begin
          end
        end
        default: stuckData_stop <= 1;
      endcase
    end
  end
  // Process: findAndInsert  process_findAndInsert_0006
  reg [6-1:0] findAndInsert_index_0;
  reg [3-1:0] findAndInsert_size_1;
  reg [1-1:0] findAndInsert_isLeaf_2;
  reg [6-1:0] findAndInsert_nextFree_3;
  reg [8-1:0] findAndInsert_Key_0_4;
  reg [1-1:0] findAndInsert_KeyCompares_0_5;
  reg [3-1:0] findAndInsert_KeyCollapse_0_6;
  reg [8-1:0] findAndInsert_Data_0_7;
  reg [8-1:0] findAndInsert_Key_1_8;
  reg [1-1:0] findAndInsert_KeyCompares_1_9;
  reg [3-1:0] findAndInsert_KeyCollapse_1_10;
  reg [8-1:0] findAndInsert_Data_1_11;
  reg [8-1:0] findAndInsert_Key_2_12;
  reg [1-1:0] findAndInsert_KeyCompares_2_13;
  reg [3-1:0] findAndInsert_KeyCollapse_2_14;
  reg [8-1:0] findAndInsert_Data_2_15;
  reg [8-1:0] findAndInsert_Key_3_16;
  reg [1-1:0] findAndInsert_KeyCompares_3_17;
  reg [3-1:0] findAndInsert_KeyCollapse_3_18;
  reg [8-1:0] findAndInsert_Data_3_19;
  reg [5-1:0] findAndInsert_stuckKeys_1_index_20;
  reg [5-1:0] findAndInsert_stuckKeys_2_index_21;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_22;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_23;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_24;
  reg [8-1:0] findAndInsert_stuckKeys_2_value_25;
  reg [5-1:0] findAndInsert_stuckData_3_index_26;
  reg [5-1:0] findAndInsert_stuckData_4_index_27;
  reg [8-1:0] findAndInsert_stuckData_4_value_28;
  reg [8-1:0] findAndInsert_stuckData_4_value_29;
  reg [8-1:0] findAndInsert_stuckData_4_value_30;
  reg [8-1:0] findAndInsert_stuckData_4_value_31;
  reg [5-1:0] findAndInsert_stuckSize_5_index_32;
  reg [5-1:0] findAndInsert_stuckSize_6_index_33;
  reg [3-1:0] findAndInsert_stuckSize_6_value_34;
  reg [5-1:0] findAndInsert_stuckIsLeaf_7_index_35;
  reg [5-1:0] findAndInsert_stuckIsLeaf_8_index_36;
  reg [1-1:0] findAndInsert_stuckIsLeaf_8_value_37;
  reg [1-1:0] findAndInsert_Found_38;
  reg [8-1:0] findAndInsert_Key_39;
  reg [8-1:0] findAndInsert_FoundKey_40;
  reg [8-1:0] findAndInsert_Data_41;
  reg [6-1:0] findAndInsert_BtreeIndex_42;
  reg [3-1:0] findAndInsert_StuckIndex_43;
  reg [1-1:0] findAndInsert_MergeSuccess_44;
  reg [6-1:0] findAndInsert_i_45;
  reg [3-1:0] findAndInsert_j_46;
  reg [6-1:0] findAndInsert_index_47;
  reg [3-1:0] findAndInsert_size_48;
  reg [1-1:0] findAndInsert_isLeaf_49;
  reg [6-1:0] findAndInsert_nextFree_50;
  reg [8-1:0] findAndInsert_Key_0_51;
  reg [1-1:0] findAndInsert_KeyCompares_0_52;
  reg [3-1:0] findAndInsert_KeyCollapse_0_53;
  reg [8-1:0] findAndInsert_Data_0_54;
  reg [8-1:0] findAndInsert_Key_1_55;
  reg [1-1:0] findAndInsert_KeyCompares_1_56;
  reg [3-1:0] findAndInsert_KeyCollapse_1_57;
  reg [8-1:0] findAndInsert_Data_1_58;
  reg [8-1:0] findAndInsert_Key_2_59;
  reg [1-1:0] findAndInsert_KeyCompares_2_60;
  reg [3-1:0] findAndInsert_KeyCollapse_2_61;
  reg [8-1:0] findAndInsert_Data_2_62;
  reg [8-1:0] findAndInsert_Key_3_63;
  reg [1-1:0] findAndInsert_KeyCompares_3_64;
  reg [3-1:0] findAndInsert_KeyCollapse_3_65;
  reg [8-1:0] findAndInsert_Data_3_66;
  reg [1-1:0] findAndInsert_Found_67;
  reg [8-1:0] findAndInsert_Key_68;
  reg [8-1:0] findAndInsert_FoundKey_69;
  reg [8-1:0] findAndInsert_Data_70;
  reg [6-1:0] findAndInsert_BtreeIndex_71;
  reg [3-1:0] findAndInsert_StuckIndex_72;
  reg [1-1:0] findAndInsert_MergeSuccess_73;
  reg [6-1:0] findAndInsert_index_74;
  reg [3-1:0] findAndInsert_size_75;
  reg [1-1:0] findAndInsert_isLeaf_76;
  reg [6-1:0] findAndInsert_nextFree_77;
  reg [8-1:0] findAndInsert_Key_0_78;
  reg [1-1:0] findAndInsert_KeyCompares_0_79;
  reg [3-1:0] findAndInsert_KeyCollapse_0_80;
  reg [8-1:0] findAndInsert_Data_0_81;
  reg [8-1:0] findAndInsert_Key_1_82;
  reg [1-1:0] findAndInsert_KeyCompares_1_83;
  reg [3-1:0] findAndInsert_KeyCollapse_1_84;
  reg [8-1:0] findAndInsert_Data_1_85;
  reg [8-1:0] findAndInsert_Key_2_86;
  reg [1-1:0] findAndInsert_KeyCompares_2_87;
  reg [3-1:0] findAndInsert_KeyCollapse_2_88;
  reg [8-1:0] findAndInsert_Data_2_89;
  reg [8-1:0] findAndInsert_Key_3_90;
  reg [1-1:0] findAndInsert_KeyCompares_3_91;
  reg [3-1:0] findAndInsert_KeyCollapse_3_92;
  reg [8-1:0] findAndInsert_Data_3_93;
  reg [1-1:0] findAndInsert_Found_94;
  reg [8-1:0] findAndInsert_Key_95;
  reg [8-1:0] findAndInsert_FoundKey_96;
  reg [8-1:0] findAndInsert_Data_97;
  reg [6-1:0] findAndInsert_BtreeIndex_98;
  reg [3-1:0] findAndInsert_StuckIndex_99;
  reg [1-1:0] findAndInsert_MergeSuccess_100;
  reg [6-1:0] findAndInsert_index_101;
  reg [3-1:0] findAndInsert_size_102;
  reg [1-1:0] findAndInsert_isLeaf_103;
  reg [6-1:0] findAndInsert_nextFree_104;
  reg [8-1:0] findAndInsert_Key_0_105;
  reg [1-1:0] findAndInsert_KeyCompares_0_106;
  reg [3-1:0] findAndInsert_KeyCollapse_0_107;
  reg [8-1:0] findAndInsert_Data_0_108;
  reg [8-1:0] findAndInsert_Key_1_109;
  reg [1-1:0] findAndInsert_KeyCompares_1_110;
  reg [3-1:0] findAndInsert_KeyCollapse_1_111;
  reg [8-1:0] findAndInsert_Data_1_112;
  reg [8-1:0] findAndInsert_Key_2_113;
  reg [1-1:0] findAndInsert_KeyCompares_2_114;
  reg [3-1:0] findAndInsert_KeyCollapse_2_115;
  reg [8-1:0] findAndInsert_Data_2_116;
  reg [8-1:0] findAndInsert_Key_3_117;
  reg [1-1:0] findAndInsert_KeyCompares_3_118;
  reg [3-1:0] findAndInsert_KeyCollapse_3_119;
  reg [8-1:0] findAndInsert_Data_3_120;
  reg [1-1:0] findAndInsert_Found_121;
  reg [8-1:0] findAndInsert_Key_122;
  reg [8-1:0] findAndInsert_FoundKey_123;
  reg [8-1:0] findAndInsert_Data_124;
  reg [6-1:0] findAndInsert_BtreeIndex_125;
  reg [3-1:0] findAndInsert_StuckIndex_126;
  reg [1-1:0] findAndInsert_MergeSuccess_127;
  reg [6-1:0] findAndInsert_index_128;
  reg [3-1:0] findAndInsert_size_129;
  reg [1-1:0] findAndInsert_isLeaf_130;
  reg [6-1:0] findAndInsert_nextFree_131;
  reg [8-1:0] findAndInsert_Key_0_132;
  reg [1-1:0] findAndInsert_KeyCompares_0_133;
  reg [3-1:0] findAndInsert_KeyCollapse_0_134;
  reg [8-1:0] findAndInsert_Data_0_135;
  reg [8-1:0] findAndInsert_Key_1_136;
  reg [1-1:0] findAndInsert_KeyCompares_1_137;
  reg [3-1:0] findAndInsert_KeyCollapse_1_138;
  reg [8-1:0] findAndInsert_Data_1_139;
  reg [8-1:0] findAndInsert_Key_2_140;
  reg [1-1:0] findAndInsert_KeyCompares_2_141;
  reg [3-1:0] findAndInsert_KeyCollapse_2_142;
  reg [8-1:0] findAndInsert_Data_2_143;
  reg [8-1:0] findAndInsert_Key_3_144;
  reg [1-1:0] findAndInsert_KeyCompares_3_145;
  reg [3-1:0] findAndInsert_KeyCollapse_3_146;
  reg [8-1:0] findAndInsert_Data_3_147;
  reg [1-1:0] findAndInsert_Found_148;
  reg [8-1:0] findAndInsert_Key_149;
  reg [8-1:0] findAndInsert_FoundKey_150;
  reg [8-1:0] findAndInsert_Data_151;
  reg [6-1:0] findAndInsert_BtreeIndex_152;
  reg [3-1:0] findAndInsert_StuckIndex_153;
  reg [1-1:0] findAndInsert_MergeSuccess_154;
  reg [8-1:0] findAndInsert_childKey_155;
  reg [6-1:0] findAndInsert_childData_156;
  reg [6-1:0] findAndInsert_indexLeft_157;
  reg [6-1:0] findAndInsert_indexRight_158;
  reg [8-1:0] findAndInsert_midKey_159;
  reg [5-1:0] findAndInsert_freeNext_9_index_160;
  reg [5-1:0] findAndInsert_freeNext_10_index_161;
  reg [6-1:0] findAndInsert_freeNext_10_value_162;
  reg [5-1:0] findAndInsert_stuckIsFree_11_index_163;
  reg [1-1:0] findAndInsert_stuckIsFree_11_value_164;
  reg [6-1:0] findAndInsert_root_165;
  reg [6-1:0] findAndInsert_next_166;
  reg [1-1:0] findAndInsert_isLeaf_167;
  reg [1-1:0] findAndInsert_isFree_168;
  reg [6-1:0] findAndInsert_index_169;
  reg [3-1:0] findAndInsert_size_170;
  reg [1-1:0] findAndInsert_isLeaf_171;
  reg [6-1:0] findAndInsert_nextFree_172;
  reg [8-1:0] findAndInsert_Key_0_173;
  reg [1-1:0] findAndInsert_KeyCompares_0_174;
  reg [3-1:0] findAndInsert_KeyCollapse_0_175;
  reg [8-1:0] findAndInsert_Data_0_176;
  reg [8-1:0] findAndInsert_Key_1_177;
  reg [1-1:0] findAndInsert_KeyCompares_1_178;
  reg [3-1:0] findAndInsert_KeyCollapse_1_179;
  reg [8-1:0] findAndInsert_Data_1_180;
  reg [8-1:0] findAndInsert_Key_2_181;
  reg [1-1:0] findAndInsert_KeyCompares_2_182;
  reg [3-1:0] findAndInsert_KeyCollapse_2_183;
  reg [8-1:0] findAndInsert_Data_2_184;
  reg [8-1:0] findAndInsert_Key_3_185;
  reg [1-1:0] findAndInsert_KeyCompares_3_186;
  reg [3-1:0] findAndInsert_KeyCollapse_3_187;
  reg [8-1:0] findAndInsert_Data_3_188;
  reg [1-1:0] findAndInsert_Found_189;
  reg [8-1:0] findAndInsert_Key_190;
  reg [8-1:0] findAndInsert_FoundKey_191;
  reg [8-1:0] findAndInsert_Data_192;
  reg [6-1:0] findAndInsert_BtreeIndex_193;
  reg [3-1:0] findAndInsert_StuckIndex_194;
  reg [1-1:0] findAndInsert_MergeSuccess_195;
  reg [6-1:0] findAndInsert_index_196;
  reg [3-1:0] findAndInsert_size_197;
  reg [1-1:0] findAndInsert_isLeaf_198;
  reg [6-1:0] findAndInsert_nextFree_199;
  reg [8-1:0] findAndInsert_Key_0_200;
  reg [1-1:0] findAndInsert_KeyCompares_0_201;
  reg [3-1:0] findAndInsert_KeyCollapse_0_202;
  reg [8-1:0] findAndInsert_Data_0_203;
  reg [8-1:0] findAndInsert_Key_1_204;
  reg [1-1:0] findAndInsert_KeyCompares_1_205;
  reg [3-1:0] findAndInsert_KeyCollapse_1_206;
  reg [8-1:0] findAndInsert_Data_1_207;
  reg [8-1:0] findAndInsert_Key_2_208;
  reg [1-1:0] findAndInsert_KeyCompares_2_209;
  reg [3-1:0] findAndInsert_KeyCollapse_2_210;
  reg [8-1:0] findAndInsert_Data_2_211;
  reg [8-1:0] findAndInsert_Key_3_212;
  reg [1-1:0] findAndInsert_KeyCompares_3_213;
  reg [3-1:0] findAndInsert_KeyCollapse_3_214;
  reg [8-1:0] findAndInsert_Data_3_215;
  reg [1-1:0] findAndInsert_Found_216;
  reg [8-1:0] findAndInsert_Key_217;
  reg [8-1:0] findAndInsert_FoundKey_218;
  reg [8-1:0] findAndInsert_Data_219;
  reg [6-1:0] findAndInsert_BtreeIndex_220;
  reg [3-1:0] findAndInsert_StuckIndex_221;
  reg [1-1:0] findAndInsert_MergeSuccess_222;
  reg [8-1:0] findAndInsert_childKey_223;
  reg [3-1:0] findAndInsert_size_224;
  reg [6-1:0] findAndInsert_childData_225;
  reg [6-1:0] findAndInsert_indexLeft_226;
  reg [6-1:0] findAndInsert_indexRight_227;
  reg [8-1:0] findAndInsert_midKey_228;
  reg [1-1:0] findAndInsert_success_229;
  reg [1-1:0] findAndInsert_test_230;
  reg [6-1:0] findAndInsert_next_231;
  reg [6-1:0] findAndInsert_root_232;
  reg [1-1:0] findAndInsert_isFree_233;
  integer findAndInsert_pc;
  integer findAndInsert_stop;
  integer findAndInsert_returnCode;
  integer findAndInsert_memory_index;
  always @ (posedge clock) begin
    if (step < 0) begin
      findAndInsert_pc <= 0;
      findAndInsert_stop <= 0;
      findAndInsert_returnCode <= 0;
      findAndInsert_index_0 <= 0;
      findAndInsert_size_1 <= 0;
      findAndInsert_isLeaf_2 <= 0;
      findAndInsert_nextFree_3 <= 0;
      findAndInsert_Key_0_4 <= 0;
      findAndInsert_KeyCompares_0_5 <= 0;
      findAndInsert_KeyCollapse_0_6 <= 0;
      findAndInsert_Data_0_7 <= 0;
      findAndInsert_Key_1_8 <= 0;
      findAndInsert_KeyCompares_1_9 <= 0;
      findAndInsert_KeyCollapse_1_10 <= 0;
      findAndInsert_Data_1_11 <= 0;
      findAndInsert_Key_2_12 <= 0;
      findAndInsert_KeyCompares_2_13 <= 0;
      findAndInsert_KeyCollapse_2_14 <= 0;
      findAndInsert_Data_2_15 <= 0;
      findAndInsert_Key_3_16 <= 0;
      findAndInsert_KeyCompares_3_17 <= 0;
      findAndInsert_KeyCollapse_3_18 <= 0;
      findAndInsert_Data_3_19 <= 0;
      findAndInsert_stuckKeys_1_index_20 <= 0;
      findAndInsert_stuckKeys_2_index_21 <= 0;
      findAndInsert_stuckKeys_2_value_22 <= 0;
      findAndInsert_stuckKeys_2_value_23 <= 0;
      findAndInsert_stuckKeys_2_value_24 <= 0;
      findAndInsert_stuckKeys_2_value_25 <= 0;
      findAndInsert_stuckData_3_index_26 <= 0;
      findAndInsert_stuckData_4_index_27 <= 0;
      findAndInsert_stuckData_4_value_28 <= 0;
      findAndInsert_stuckData_4_value_29 <= 0;
      findAndInsert_stuckData_4_value_30 <= 0;
      findAndInsert_stuckData_4_value_31 <= 0;
      findAndInsert_stuckSize_5_index_32 <= 0;
      findAndInsert_stuckSize_6_index_33 <= 0;
      findAndInsert_stuckSize_6_value_34 <= 0;
      findAndInsert_stuckIsLeaf_7_index_35 <= 0;
      findAndInsert_stuckIsLeaf_8_index_36 <= 0;
      findAndInsert_stuckIsLeaf_8_value_37 <= 0;
      findAndInsert_Found_38 <= 0;
      findAndInsert_Key_39 <= 0;
      findAndInsert_FoundKey_40 <= 0;
      findAndInsert_Data_41 <= 0;
      findAndInsert_BtreeIndex_42 <= 0;
      findAndInsert_StuckIndex_43 <= 0;
      findAndInsert_MergeSuccess_44 <= 0;
      findAndInsert_i_45 <= 0;
      findAndInsert_j_46 <= 0;
      findAndInsert_index_47 <= 0;
      findAndInsert_size_48 <= 0;
      findAndInsert_isLeaf_49 <= 0;
      findAndInsert_nextFree_50 <= 0;
      findAndInsert_Key_0_51 <= 0;
      findAndInsert_KeyCompares_0_52 <= 0;
      findAndInsert_KeyCollapse_0_53 <= 0;
      findAndInsert_Data_0_54 <= 0;
      findAndInsert_Key_1_55 <= 0;
      findAndInsert_KeyCompares_1_56 <= 0;
      findAndInsert_KeyCollapse_1_57 <= 0;
      findAndInsert_Data_1_58 <= 0;
      findAndInsert_Key_2_59 <= 0;
      findAndInsert_KeyCompares_2_60 <= 0;
      findAndInsert_KeyCollapse_2_61 <= 0;
      findAndInsert_Data_2_62 <= 0;
      findAndInsert_Key_3_63 <= 0;
      findAndInsert_KeyCompares_3_64 <= 0;
      findAndInsert_KeyCollapse_3_65 <= 0;
      findAndInsert_Data_3_66 <= 0;
      findAndInsert_Found_67 <= 0;
      findAndInsert_Key_68 <= 0;
      findAndInsert_FoundKey_69 <= 0;
      findAndInsert_Data_70 <= 0;
      findAndInsert_BtreeIndex_71 <= 0;
      findAndInsert_StuckIndex_72 <= 0;
      findAndInsert_MergeSuccess_73 <= 0;
      findAndInsert_index_74 <= 0;
      findAndInsert_size_75 <= 0;
      findAndInsert_isLeaf_76 <= 0;
      findAndInsert_nextFree_77 <= 0;
      findAndInsert_Key_0_78 <= 0;
      findAndInsert_KeyCompares_0_79 <= 0;
      findAndInsert_KeyCollapse_0_80 <= 0;
      findAndInsert_Data_0_81 <= 0;
      findAndInsert_Key_1_82 <= 0;
      findAndInsert_KeyCompares_1_83 <= 0;
      findAndInsert_KeyCollapse_1_84 <= 0;
      findAndInsert_Data_1_85 <= 0;
      findAndInsert_Key_2_86 <= 0;
      findAndInsert_KeyCompares_2_87 <= 0;
      findAndInsert_KeyCollapse_2_88 <= 0;
      findAndInsert_Data_2_89 <= 0;
      findAndInsert_Key_3_90 <= 0;
      findAndInsert_KeyCompares_3_91 <= 0;
      findAndInsert_KeyCollapse_3_92 <= 0;
      findAndInsert_Data_3_93 <= 0;
      findAndInsert_Found_94 <= 0;
      findAndInsert_Key_95 <= 0;
      findAndInsert_FoundKey_96 <= 0;
      findAndInsert_Data_97 <= 0;
      findAndInsert_BtreeIndex_98 <= 0;
      findAndInsert_StuckIndex_99 <= 0;
      findAndInsert_MergeSuccess_100 <= 0;
      findAndInsert_index_101 <= 0;
      findAndInsert_size_102 <= 0;
      findAndInsert_isLeaf_103 <= 0;
      findAndInsert_nextFree_104 <= 0;
      findAndInsert_Key_0_105 <= 0;
      findAndInsert_KeyCompares_0_106 <= 0;
      findAndInsert_KeyCollapse_0_107 <= 0;
      findAndInsert_Data_0_108 <= 0;
      findAndInsert_Key_1_109 <= 0;
      findAndInsert_KeyCompares_1_110 <= 0;
      findAndInsert_KeyCollapse_1_111 <= 0;
      findAndInsert_Data_1_112 <= 0;
      findAndInsert_Key_2_113 <= 0;
      findAndInsert_KeyCompares_2_114 <= 0;
      findAndInsert_KeyCollapse_2_115 <= 0;
      findAndInsert_Data_2_116 <= 0;
      findAndInsert_Key_3_117 <= 0;
      findAndInsert_KeyCompares_3_118 <= 0;
      findAndInsert_KeyCollapse_3_119 <= 0;
      findAndInsert_Data_3_120 <= 0;
      findAndInsert_Found_121 <= 0;
      findAndInsert_Key_122 <= 0;
      findAndInsert_FoundKey_123 <= 0;
      findAndInsert_Data_124 <= 0;
      findAndInsert_BtreeIndex_125 <= 0;
      findAndInsert_StuckIndex_126 <= 0;
      findAndInsert_MergeSuccess_127 <= 0;
      findAndInsert_index_128 <= 0;
      findAndInsert_size_129 <= 0;
      findAndInsert_isLeaf_130 <= 0;
      findAndInsert_nextFree_131 <= 0;
      findAndInsert_Key_0_132 <= 0;
      findAndInsert_KeyCompares_0_133 <= 0;
      findAndInsert_KeyCollapse_0_134 <= 0;
      findAndInsert_Data_0_135 <= 0;
      findAndInsert_Key_1_136 <= 0;
      findAndInsert_KeyCompares_1_137 <= 0;
      findAndInsert_KeyCollapse_1_138 <= 0;
      findAndInsert_Data_1_139 <= 0;
      findAndInsert_Key_2_140 <= 0;
      findAndInsert_KeyCompares_2_141 <= 0;
      findAndInsert_KeyCollapse_2_142 <= 0;
      findAndInsert_Data_2_143 <= 0;
      findAndInsert_Key_3_144 <= 0;
      findAndInsert_KeyCompares_3_145 <= 0;
      findAndInsert_KeyCollapse_3_146 <= 0;
      findAndInsert_Data_3_147 <= 0;
      findAndInsert_Found_148 <= 0;
      findAndInsert_Key_149 <= 0;
      findAndInsert_FoundKey_150 <= 0;
      findAndInsert_Data_151 <= 0;
      findAndInsert_BtreeIndex_152 <= 0;
      findAndInsert_StuckIndex_153 <= 0;
      findAndInsert_MergeSuccess_154 <= 0;
      findAndInsert_childKey_155 <= 0;
      findAndInsert_childData_156 <= 0;
      findAndInsert_indexLeft_157 <= 0;
      findAndInsert_indexRight_158 <= 0;
      findAndInsert_midKey_159 <= 0;
      findAndInsert_freeNext_9_index_160 <= 0;
      findAndInsert_freeNext_10_index_161 <= 0;
      findAndInsert_freeNext_10_value_162 <= 0;
      findAndInsert_stuckIsFree_11_index_163 <= 0;
      findAndInsert_stuckIsFree_11_value_164 <= 0;
      findAndInsert_root_165 <= 0;
      findAndInsert_next_166 <= 0;
      findAndInsert_isLeaf_167 <= 0;
      findAndInsert_isFree_168 <= 0;
      findAndInsert_index_169 <= 0;
      findAndInsert_size_170 <= 0;
      findAndInsert_isLeaf_171 <= 0;
      findAndInsert_nextFree_172 <= 0;
      findAndInsert_Key_0_173 <= 0;
      findAndInsert_KeyCompares_0_174 <= 0;
      findAndInsert_KeyCollapse_0_175 <= 0;
      findAndInsert_Data_0_176 <= 0;
      findAndInsert_Key_1_177 <= 0;
      findAndInsert_KeyCompares_1_178 <= 0;
      findAndInsert_KeyCollapse_1_179 <= 0;
      findAndInsert_Data_1_180 <= 0;
      findAndInsert_Key_2_181 <= 0;
      findAndInsert_KeyCompares_2_182 <= 0;
      findAndInsert_KeyCollapse_2_183 <= 0;
      findAndInsert_Data_2_184 <= 0;
      findAndInsert_Key_3_185 <= 0;
      findAndInsert_KeyCompares_3_186 <= 0;
      findAndInsert_KeyCollapse_3_187 <= 0;
      findAndInsert_Data_3_188 <= 0;
      findAndInsert_Found_189 <= 0;
      findAndInsert_Key_190 <= 0;
      findAndInsert_FoundKey_191 <= 0;
      findAndInsert_Data_192 <= 0;
      findAndInsert_BtreeIndex_193 <= 0;
      findAndInsert_StuckIndex_194 <= 0;
      findAndInsert_MergeSuccess_195 <= 0;
      findAndInsert_index_196 <= 0;
      findAndInsert_size_197 <= 0;
      findAndInsert_isLeaf_198 <= 0;
      findAndInsert_nextFree_199 <= 0;
      findAndInsert_Key_0_200 <= 0;
      findAndInsert_KeyCompares_0_201 <= 0;
      findAndInsert_KeyCollapse_0_202 <= 0;
      findAndInsert_Data_0_203 <= 0;
      findAndInsert_Key_1_204 <= 0;
      findAndInsert_KeyCompares_1_205 <= 0;
      findAndInsert_KeyCollapse_1_206 <= 0;
      findAndInsert_Data_1_207 <= 0;
      findAndInsert_Key_2_208 <= 0;
      findAndInsert_KeyCompares_2_209 <= 0;
      findAndInsert_KeyCollapse_2_210 <= 0;
      findAndInsert_Data_2_211 <= 0;
      findAndInsert_Key_3_212 <= 0;
      findAndInsert_KeyCompares_3_213 <= 0;
      findAndInsert_KeyCollapse_3_214 <= 0;
      findAndInsert_Data_3_215 <= 0;
      findAndInsert_Found_216 <= 0;
      findAndInsert_Key_217 <= 0;
      findAndInsert_FoundKey_218 <= 0;
      findAndInsert_Data_219 <= 0;
      findAndInsert_BtreeIndex_220 <= 0;
      findAndInsert_StuckIndex_221 <= 0;
      findAndInsert_MergeSuccess_222 <= 0;
      findAndInsert_childKey_223 <= 0;
      findAndInsert_size_224 <= 0;
      findAndInsert_childData_225 <= 0;
      findAndInsert_indexLeft_226 <= 0;
      findAndInsert_indexRight_227 <= 0;
      findAndInsert_midKey_228 <= 0;
      findAndInsert_success_229 <= 0;
      findAndInsert_test_230 <= 0;
      findAndInsert_next_231 <= 0;
      findAndInsert_root_232 <= 0;
      findAndInsert_isFree_233 <= 0;
      stuckIsLeaf_7_requestedAt <= -1;
      stuckIsLeaf_8_requestedAt <= -1;
      stuckIsFree_11_requestedAt <= -1;
      freeNext_9_requestedAt <= -1;
      freeNext_10_requestedAt <= -1;
      stuckSize_5_requestedAt <= -1;
      stuckSize_6_requestedAt <= -1;
      stuckKeys_1_requestedAt <= -1;
      stuckKeys_2_requestedAt <= -1;
      stuckData_3_requestedAt <= -1;
      stuckData_4_requestedAt <= -1;
    end
    else if (processCurrent == 6) begin
      case(findAndInsert_pc)
        0: begin
          findAndInsert_i_45 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0676:<init>|  Chip.java:0675:RegisterSet|  Btree.java:4580:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        1: begin
          findAndInsert_index_0 <= findAndInsert_i_45;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        2: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_0;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_0;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_0;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_0;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        3: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        4: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        5: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        6: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        7: begin
          findAndInsert_size_1 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_2 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_4 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_7 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_8 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_11 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_12 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_15 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_16 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_19 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:4581:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        8: begin
          if (findAndInsert_i_45 == 0 && findAndInsert_size_1 > 1) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          else begin
            if (findAndInsert_i_45 == 0 || findAndInsert_size_1 < 1) begin
              findAndInsert_pc <= 53;
            end
            else begin
              findAndInsert_pc <= findAndInsert_pc + 1;
            end
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1768:<init>|  Btree.java:1767:mergePermitted|  Btree.java:2183:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        9: begin
          findAndInsert_success_229 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:2184:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        10: begin
          findAndInsert_size_224 <= findAndInsert_size_1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:2185:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        11: begin
          case (findAndInsert_size_224)
            1: begin
              findAndInsert_indexLeft_226 <= findAndInsert_Data_0_7;
              findAndInsert_indexRight_227 <= findAndInsert_Data_1_11;
            end
            2: begin
              findAndInsert_indexLeft_226 <= findAndInsert_Data_1_11;
              findAndInsert_indexRight_227 <= findAndInsert_Data_2_15;
            end
            3: begin
              findAndInsert_indexLeft_226 <= findAndInsert_Data_2_15;
              findAndInsert_indexRight_227 <= findAndInsert_Data_3_19;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2188:<init>|  Btree.java:2187:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        12: begin
          findAndInsert_index_169 <= findAndInsert_indexLeft_226;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        13: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_169;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_169;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_169;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_169;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        14: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        15: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        16: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        17: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        18: begin
          findAndInsert_size_170 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_171 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_173 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_176 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_177 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_180 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_181 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_184 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_185 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_188 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2202:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        19: begin
          findAndInsert_index_196 <= findAndInsert_indexRight_227;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0697:<init>|  Chip.java:0696:Copy|  Btree.java:0261:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        20: begin
          findAndInsert_stuckSize_5_index_32 <= findAndInsert_index_196;
          stuckSize_5_requestedAt <= step;
          stuckSize_5_finishedAt <= -1;
          findAndInsert_stuckIsLeaf_7_index_35 <= findAndInsert_index_196;
          stuckIsLeaf_7_requestedAt <= step;
          stuckIsLeaf_7_finishedAt <= -1;
          findAndInsert_stuckKeys_1_index_20 <= findAndInsert_index_196;
          stuckKeys_1_requestedAt <= step;
          stuckKeys_1_finishedAt <= -1;
          findAndInsert_stuckData_3_index_26 <= findAndInsert_index_196;
          stuckData_3_requestedAt <= step;
          stuckData_3_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0272:<init>|  Btree.java:0271:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        21: begin
          if ((stuckSize_5_requestedAt < stuckSize_5_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0285:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        22: begin
          if ((stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0286:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        23: begin
          if ((stuckKeys_1_requestedAt < stuckKeys_1_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0288:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        24: begin
          if ((stuckData_3_requestedAt < stuckData_3_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0289:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        25: begin
          findAndInsert_size_197 <= stuckSize_stuckSize_5_result_0;
          findAndInsert_isLeaf_198 <= stuckIsLeaf_stuckIsLeaf_7_result_0;
          findAndInsert_Key_0_200 <= stuckKeys_stuckKeys_1_result_0;
          findAndInsert_Data_0_203 <= stuckData_stuckData_3_result_0;
          findAndInsert_Key_1_204 <= stuckKeys_stuckKeys_1_result_1;
          findAndInsert_Data_1_207 <= stuckData_stuckData_3_result_1;
          findAndInsert_Key_2_208 <= stuckKeys_stuckKeys_1_result_2;
          findAndInsert_Data_2_211 <= stuckData_stuckData_3_result_2;
          findAndInsert_Key_3_212 <= stuckKeys_stuckKeys_1_result_3;
          findAndInsert_Data_3_215 <= stuckData_stuckData_3_result_3;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0292:<init>|  Btree.java:0291:stuckGet|  Btree.java:0262:stuckGet|  Btree.java:2203:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        26: begin
          if (findAndInsert_isLeaf_171 == 0) begin
            findAndInsert_pc <= 28;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        27: begin
          findAndInsert_pc <= 53;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        28: begin
          if (findAndInsert_isLeaf_198 == 0) begin
            findAndInsert_pc <= 30;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Btree.java:1394:<init>|  Btree.java:1393:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        29: begin
          findAndInsert_pc <= 53;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0571:<init>|  Chip.java:0570:GOto|  Btree.java:1410:code|  Chip.java:0530:<init>|  Btree.java:1391:<init>|  Btree.java:1390:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        30: begin
          case (findAndInsert_size_1)
            1: begin
              findAndInsert_Key_39 <= findAndInsert_Key_0_4;
              findAndInsert_Data_41 <= findAndInsert_Data_0_7;
            end
            2: begin
              findAndInsert_Key_39 <= findAndInsert_Key_1_8;
              findAndInsert_Data_41 <= findAndInsert_Data_1_11;
            end
            3: begin
              findAndInsert_Key_39 <= findAndInsert_Key_2_12;
              findAndInsert_Data_41 <= findAndInsert_Data_2_15;
            end
            4: begin
              findAndInsert_Key_39 <= findAndInsert_Key_3_16;
              findAndInsert_Data_41 <= findAndInsert_Data_3_19;
            end
          endcase
          findAndInsert_size_1 <= findAndInsert_size_1-1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0452:<init>|  Btree.java:0451:Pop|  Btree.java:2209:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        31: begin
          findAndInsert_MergeSuccess_195 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:1286:mergeButOne|  Btree.java:2210:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        32: begin
          case (findAndInsert_size_170)
            0: begin
              case (findAndInsert_size_197)
                0: begin
                  findAndInsert_Key_0_173 <= findAndInsert_Key_39;
                  findAndInsert_Data_1_180 <= findAndInsert_Data_0_203;
                  findAndInsert_size_170 <= findAndInsert_size_170 + 1;
                  findAndInsert_MergeSuccess_195 <= 1;
                end
                1: begin
                  findAndInsert_Key_0_173 <= findAndInsert_Key_39;
                  findAndInsert_Key_1_177 <= findAndInsert_Key_0_200;
                  findAndInsert_Data_1_180 <= findAndInsert_Data_0_203;
                  findAndInsert_Data_2_184 <= findAndInsert_Data_1_207;
                  findAndInsert_size_170 <= findAndInsert_size_170 + 2;
                  findAndInsert_MergeSuccess_195 <= 1;
                end
                2: begin
                  findAndInsert_Key_0_173 <= findAndInsert_Key_39;
                  findAndInsert_Key_1_177 <= findAndInsert_Key_0_200;
                  findAndInsert_Data_1_180 <= findAndInsert_Data_0_203;
                  findAndInsert_Key_2_181 <= findAndInsert_Key_1_204;
                  findAndInsert_Data_2_184 <= findAndInsert_Data_1_207;
                  findAndInsert_Data_3_188 <= findAndInsert_Data_2_211;
                  findAndInsert_size_170 <= findAndInsert_size_170 + 3;
                  findAndInsert_MergeSuccess_195 <= 1;
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            1: begin
              case (findAndInsert_size_197)
                0: begin
                  findAndInsert_Key_1_177 <= findAndInsert_Key_39;
                  findAndInsert_Data_2_184 <= findAndInsert_Data_0_203;
                  findAndInsert_size_170 <= findAndInsert_size_170 + 1;
                  findAndInsert_MergeSuccess_195 <= 1;
                end
                1: begin
                  findAndInsert_Key_1_177 <= findAndInsert_Key_39;
                  findAndInsert_Key_2_181 <= findAndInsert_Key_0_200;
                  findAndInsert_Data_2_184 <= findAndInsert_Data_0_203;
                  findAndInsert_Data_3_188 <= findAndInsert_Data_1_207;
                  findAndInsert_size_170 <= findAndInsert_size_170 + 2;
                  findAndInsert_MergeSuccess_195 <= 1;
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            2: begin
              case (findAndInsert_size_197)
                0: begin
                  findAndInsert_Key_2_181 <= findAndInsert_Key_39;
                  findAndInsert_Data_3_188 <= findAndInsert_Data_0_203;
                  findAndInsert_size_170 <= findAndInsert_size_170 + 1;
                  findAndInsert_MergeSuccess_195 <= 1;
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            3: begin
              case (findAndInsert_size_197)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
            4: begin
              case (findAndInsert_size_197)
                0: begin
                end
                1: begin
                end
                2: begin
                end
                3: begin
                end
                4: begin
                end
              endcase
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:1288:<init>|  Btree.java:1287:mergeButOne|  Btree.java:2210:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        33: begin
          if (findAndInsert_MergeSuccess_195 == 0) begin
            findAndInsert_pc <= 53;
          end
          else begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0603:<init>|  Chip.java:0602:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        34: begin
          findAndInsert_success_229 <= 1;
          case (findAndInsert_size_1)
            0: begin
              findAndInsert_Key_0_4 <= findAndInsert_Key_39;
              findAndInsert_Data_0_7 <= findAndInsert_indexLeft_226;
            end
            1: begin
              findAndInsert_Key_1_8 <= findAndInsert_Key_39;
              findAndInsert_Data_1_11 <= findAndInsert_indexLeft_226;
            end
            2: begin
              findAndInsert_Key_2_12 <= findAndInsert_Key_39;
              findAndInsert_Data_2_15 <= findAndInsert_indexLeft_226;
            end
            3: begin
              findAndInsert_Key_3_16 <= findAndInsert_Key_39;
              findAndInsert_Data_3_19 <= findAndInsert_indexLeft_226;
            end
          endcase
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:2214:<init>|  Btree.java:2213:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        35: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_169;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_170;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_169;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_173;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_177;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_181;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_185;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_169;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_176;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_180;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_184;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_188;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        36: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        37: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        38: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2224:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        39: begin
          findAndInsert_stuckSize_6_index_33 <= findAndInsert_index_0;
          findAndInsert_stuckSize_6_value_34 <= findAndInsert_size_1;
          stuckSize_6_requestedAt <= step;
          stuckSize_6_finishedAt <= -1;
          findAndInsert_stuckKeys_2_index_21 <= findAndInsert_index_0;
          findAndInsert_stuckKeys_2_value_22 <= findAndInsert_Key_0_4;
          findAndInsert_stuckKeys_2_value_23 <= findAndInsert_Key_1_8;
          findAndInsert_stuckKeys_2_value_24 <= findAndInsert_Key_2_12;
          findAndInsert_stuckKeys_2_value_25 <= findAndInsert_Key_3_16;
          stuckKeys_2_requestedAt <= step;
          stuckKeys_2_finishedAt <= -1;
          findAndInsert_stuckData_4_index_27 <= findAndInsert_index_0;
          findAndInsert_stuckData_4_value_28 <= findAndInsert_Data_0_7;
          findAndInsert_stuckData_4_value_29 <= findAndInsert_Data_1_11;
          findAndInsert_stuckData_4_value_30 <= findAndInsert_Data_2_15;
          findAndInsert_stuckData_4_value_31 <= findAndInsert_Data_3_19;
          stuckData_4_requestedAt <= step;
          stuckData_4_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0313:<init>|  Btree.java:0312:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        40: begin
          if ((stuckSize_6_requestedAt < stuckSize_6_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0327:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        41: begin
          if ((stuckKeys_2_requestedAt < stuckKeys_2_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0330:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        42: begin
          if ((stuckData_4_requestedAt < stuckData_4_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0331:stuckPut|  Btree.java:0334:stuckPut|  Btree.java:2225:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        43: begin
          findAndInsert_root_232 <= 0;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:0792:<init>|  Chip.java:0791:Zero|  Btree.java:0127:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        44: begin
          findAndInsert_freeNext_9_index_160 <= findAndInsert_root_232;
          freeNext_9_requestedAt <= step;
          freeNext_9_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1300:<init>|  Chip.java:1299:ExecuteTransaction|  Btree.java:0128:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        45: begin
          if ((freeNext_9_requestedAt < freeNext_9_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1307:<init>|  Chip.java:1306:waitResultOfTransaction|  Btree.java:0129:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        46: begin
          findAndInsert_next_231 <= freeNext_freeNext_9_result_0;
          findAndInsert_freeNext_10_index_161 <= findAndInsert_root_232;
          findAndInsert_freeNext_10_value_162 <= findAndInsert_indexRight_227;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_isFree_233 <= 1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Btree.java:0132:<init>|  Btree.java:0131:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        47: begin
          findAndInsert_stuckIsFree_11_index_163 <= findAndInsert_indexRight_227;
          findAndInsert_stuckIsFree_11_value_164 <= findAndInsert_isFree_233;
          stuckIsFree_11_requestedAt <= step;
          stuckIsFree_11_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0144:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        48: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0145:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        49: begin
          findAndInsert_freeNext_10_index_161 <= findAndInsert_indexRight_227;
          findAndInsert_freeNext_10_value_162 <= findAndInsert_next_231;
          freeNext_10_requestedAt <= step;
          freeNext_10_finishedAt <= -1;
          findAndInsert_pc <= findAndInsert_pc + 1;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0512:<init>|  Chip.java:1363:<init>|  Chip.java:1362:ExecuteTransaction|  Btree.java:0146:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        50: begin
          if ((freeNext_10_requestedAt < freeNext_10_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0147:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        51: begin
          if ((stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt)) begin
            findAndInsert_pc <= findAndInsert_pc + 1;
          end
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:1370:<init>|  Chip.java:1369:waitResultOfTransaction|  Btree.java:0148:free|  Btree.java:2226:Then|  Chip.java:0610:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        52: begin
          findAndInsert_pc <= 53;
          begin
            integer f;
            f = $fopen("verilog/trace_verilog.txt", "a");
            $fdisplay(f, "Location: Chip.java:0612:<init>|  Chip.java:0611:<init>|  Btree.java:2212:<init>|  Btree.java:2211:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2208:<init>|  Btree.java:2207:Branch|  Btree.java:1413:code|  Chip.java:0530:<init>|  Btree.java:1388:<init>|  Btree.java:1387:<init>|  Btree.java:2206:<init>|  Btree.java:2205:code|  Chip.java:0530:<init>|  Btree.java:2182:<init>|  Btree.java:2181:mergeBranchesAtTop|  Btree.java:4582:test_mergeBranchesAtTop|  Btree.java:6980:newTests|  Btree.java:6986:main|");
            $fclose(f);
          end
        end
        default: findAndInsert_stop <= 1;
      endcase
    end
  end
  task chipPrint;
    begin
      integer o;
      o = $fopen("verilog/trace_verilog.txt", "a");
      if (!o) o = $fopen("../verilog/trace_verilog.txt", "a");
      if (!o) $display("Cannot create trace folder: verilog/trace_verilog.txt");
      $fwrite(o, "Chip: %-16s step: %1d, maxSteps: %1d, running: %1d\n", "Btree", step, maxSteps, !stop);
      $fwrite(o, "  Processes:\n");

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 0, "stuckIsLeaf", 1, stuckIsLeaf_pc, stuckIsLeaf_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsLeaf_memory[0]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[1]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[2]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[3]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[4]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[5]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[6]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[7]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[8]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[9]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[10]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[11]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[12]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[13]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[14]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[15]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[16]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[17]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[18]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[19]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[20]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[21]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[22]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[23]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[24]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[25]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[26]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[27]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[28]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[29]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[30]);
      $fwrite(o, ", %2d", stuckIsLeaf_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckIsLeaf_7", stuckIsLeaf_7_requestedAt, stuckIsLeaf_7_finishedAt, stuckIsLeaf_stuckIsLeaf_7_returnCode, (stuckIsLeaf_7_requestedAt > stuckIsLeaf_7_finishedAt && stuckIsLeaf_7_requestedAt != step), (stuckIsLeaf_7_requestedAt < stuckIsLeaf_7_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsLeaf_7_index_35", findAndInsert_stuckIsLeaf_7_index_35);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckIsLeaf_stuckIsLeaf_7_result_0", stuckIsLeaf_stuckIsLeaf_7_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsLeaf_8", stuckIsLeaf_8_requestedAt, stuckIsLeaf_8_finishedAt, stuckIsLeaf_stuckIsLeaf_8_returnCode, (stuckIsLeaf_8_requestedAt > stuckIsLeaf_8_finishedAt && stuckIsLeaf_8_requestedAt != step), (stuckIsLeaf_8_requestedAt < stuckIsLeaf_8_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsLeaf_8_index_36", findAndInsert_stuckIsLeaf_8_index_36);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsLeaf_8_value_37", findAndInsert_stuckIsLeaf_8_value_37);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 1, "stuckIsFree", 1, stuckIsFree_pc, stuckIsFree_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 1, 1);
      $fwrite(o, "        %2d", stuckIsFree_memory[0]);
      $fwrite(o, ", %2d", stuckIsFree_memory[1]);
      $fwrite(o, ", %2d", stuckIsFree_memory[2]);
      $fwrite(o, ", %2d", stuckIsFree_memory[3]);
      $fwrite(o, ", %2d", stuckIsFree_memory[4]);
      $fwrite(o, ", %2d", stuckIsFree_memory[5]);
      $fwrite(o, ", %2d", stuckIsFree_memory[6]);
      $fwrite(o, ", %2d", stuckIsFree_memory[7]);
      $fwrite(o, ", %2d", stuckIsFree_memory[8]);
      $fwrite(o, ", %2d", stuckIsFree_memory[9]);
      $fwrite(o, ", %2d", stuckIsFree_memory[10]);
      $fwrite(o, ", %2d", stuckIsFree_memory[11]);
      $fwrite(o, ", %2d", stuckIsFree_memory[12]);
      $fwrite(o, ", %2d", stuckIsFree_memory[13]);
      $fwrite(o, ", %2d", stuckIsFree_memory[14]);
      $fwrite(o, ", %2d", stuckIsFree_memory[15]);
      $fwrite(o, ", %2d", stuckIsFree_memory[16]);
      $fwrite(o, ", %2d", stuckIsFree_memory[17]);
      $fwrite(o, ", %2d", stuckIsFree_memory[18]);
      $fwrite(o, ", %2d", stuckIsFree_memory[19]);
      $fwrite(o, ", %2d", stuckIsFree_memory[20]);
      $fwrite(o, ", %2d", stuckIsFree_memory[21]);
      $fwrite(o, ", %2d", stuckIsFree_memory[22]);
      $fwrite(o, ", %2d", stuckIsFree_memory[23]);
      $fwrite(o, ", %2d", stuckIsFree_memory[24]);
      $fwrite(o, ", %2d", stuckIsFree_memory[25]);
      $fwrite(o, ", %2d", stuckIsFree_memory[26]);
      $fwrite(o, ", %2d", stuckIsFree_memory[27]);
      $fwrite(o, ", %2d", stuckIsFree_memory[28]);
      $fwrite(o, ", %2d", stuckIsFree_memory[29]);
      $fwrite(o, ", %2d", stuckIsFree_memory[30]);
      $fwrite(o, ", %2d", stuckIsFree_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckIsFree_11", stuckIsFree_11_requestedAt, stuckIsFree_11_finishedAt, stuckIsFree_stuckIsFree_11_returnCode, (stuckIsFree_11_requestedAt > stuckIsFree_11_finishedAt && stuckIsFree_11_requestedAt != step), (stuckIsFree_11_requestedAt < stuckIsFree_11_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsFree_11_index_163", findAndInsert_stuckIsFree_11_index_163);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckIsFree_11_value_164", findAndInsert_stuckIsFree_11_value_164);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 2, "freeNext", 1, freeNext_pc, freeNext_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 6, 1);
      $fwrite(o, "        %2d", freeNext_memory[0]);
      $fwrite(o, ", %2d", freeNext_memory[1]);
      $fwrite(o, ", %2d", freeNext_memory[2]);
      $fwrite(o, ", %2d", freeNext_memory[3]);
      $fwrite(o, ", %2d", freeNext_memory[4]);
      $fwrite(o, ", %2d", freeNext_memory[5]);
      $fwrite(o, ", %2d", freeNext_memory[6]);
      $fwrite(o, ", %2d", freeNext_memory[7]);
      $fwrite(o, ", %2d", freeNext_memory[8]);
      $fwrite(o, ", %2d", freeNext_memory[9]);
      $fwrite(o, ", %2d", freeNext_memory[10]);
      $fwrite(o, ", %2d", freeNext_memory[11]);
      $fwrite(o, ", %2d", freeNext_memory[12]);
      $fwrite(o, ", %2d", freeNext_memory[13]);
      $fwrite(o, ", %2d", freeNext_memory[14]);
      $fwrite(o, ", %2d", freeNext_memory[15]);
      $fwrite(o, ", %2d", freeNext_memory[16]);
      $fwrite(o, ", %2d", freeNext_memory[17]);
      $fwrite(o, ", %2d", freeNext_memory[18]);
      $fwrite(o, ", %2d", freeNext_memory[19]);
      $fwrite(o, ", %2d", freeNext_memory[20]);
      $fwrite(o, ", %2d", freeNext_memory[21]);
      $fwrite(o, ", %2d", freeNext_memory[22]);
      $fwrite(o, ", %2d", freeNext_memory[23]);
      $fwrite(o, ", %2d", freeNext_memory[24]);
      $fwrite(o, ", %2d", freeNext_memory[25]);
      $fwrite(o, ", %2d", freeNext_memory[26]);
      $fwrite(o, ", %2d", freeNext_memory[27]);
      $fwrite(o, ", %2d", freeNext_memory[28]);
      $fwrite(o, ", %2d", freeNext_memory[29]);
      $fwrite(o, ", %2d", freeNext_memory[30]);
      $fwrite(o, ", %2d", freeNext_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "freeNext_9", freeNext_9_requestedAt, freeNext_9_finishedAt, freeNext_freeNext_9_returnCode, (freeNext_9_requestedAt > freeNext_9_finishedAt && freeNext_9_requestedAt != step), (freeNext_9_requestedAt < freeNext_9_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_freeNext_9_index_160", findAndInsert_freeNext_9_index_160);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "freeNext_freeNext_9_result_0", freeNext_freeNext_9_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "freeNext_10", freeNext_10_requestedAt, freeNext_10_finishedAt, freeNext_freeNext_10_returnCode, (freeNext_10_requestedAt > freeNext_10_finishedAt && freeNext_10_requestedAt != step), (freeNext_10_requestedAt < freeNext_10_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_freeNext_10_index_161", findAndInsert_freeNext_10_index_161);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_freeNext_10_value_162", findAndInsert_freeNext_10_value_162);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 3, "stuckSize", 1, stuckSize_pc, stuckSize_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 3, 1);
      $fwrite(o, "        %2d", stuckSize_memory[0]);
      $fwrite(o, ", %2d", stuckSize_memory[1]);
      $fwrite(o, ", %2d", stuckSize_memory[2]);
      $fwrite(o, ", %2d", stuckSize_memory[3]);
      $fwrite(o, ", %2d", stuckSize_memory[4]);
      $fwrite(o, ", %2d", stuckSize_memory[5]);
      $fwrite(o, ", %2d", stuckSize_memory[6]);
      $fwrite(o, ", %2d", stuckSize_memory[7]);
      $fwrite(o, ", %2d", stuckSize_memory[8]);
      $fwrite(o, ", %2d", stuckSize_memory[9]);
      $fwrite(o, ", %2d", stuckSize_memory[10]);
      $fwrite(o, ", %2d", stuckSize_memory[11]);
      $fwrite(o, ", %2d", stuckSize_memory[12]);
      $fwrite(o, ", %2d", stuckSize_memory[13]);
      $fwrite(o, ", %2d", stuckSize_memory[14]);
      $fwrite(o, ", %2d", stuckSize_memory[15]);
      $fwrite(o, ", %2d", stuckSize_memory[16]);
      $fwrite(o, ", %2d", stuckSize_memory[17]);
      $fwrite(o, ", %2d", stuckSize_memory[18]);
      $fwrite(o, ", %2d", stuckSize_memory[19]);
      $fwrite(o, ", %2d", stuckSize_memory[20]);
      $fwrite(o, ", %2d", stuckSize_memory[21]);
      $fwrite(o, ", %2d", stuckSize_memory[22]);
      $fwrite(o, ", %2d", stuckSize_memory[23]);
      $fwrite(o, ", %2d", stuckSize_memory[24]);
      $fwrite(o, ", %2d", stuckSize_memory[25]);
      $fwrite(o, ", %2d", stuckSize_memory[26]);
      $fwrite(o, ", %2d", stuckSize_memory[27]);
      $fwrite(o, ", %2d", stuckSize_memory[28]);
      $fwrite(o, ", %2d", stuckSize_memory[29]);
      $fwrite(o, ", %2d", stuckSize_memory[30]);
      $fwrite(o, ", %2d", stuckSize_memory[31]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckSize_5", stuckSize_5_requestedAt, stuckSize_5_finishedAt, stuckSize_stuckSize_5_returnCode, (stuckSize_5_requestedAt > stuckSize_5_finishedAt && stuckSize_5_requestedAt != step), (stuckSize_5_requestedAt < stuckSize_5_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckSize_5_index_32", findAndInsert_stuckSize_5_index_32);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckSize_stuckSize_5_result_0", stuckSize_stuckSize_5_result_0);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckSize_6", stuckSize_6_requestedAt, stuckSize_6_finishedAt, stuckSize_stuckSize_6_returnCode, (stuckSize_6_requestedAt > stuckSize_6_finishedAt && stuckSize_6_requestedAt != step), (stuckSize_6_requestedAt < stuckSize_6_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckSize_6_index_33", findAndInsert_stuckSize_6_index_33);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckSize_6_value_34", findAndInsert_stuckSize_6_value_34);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 4, "stuckKeys", 1, stuckKeys_pc, stuckKeys_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckKeys_memory[0]);
      $fwrite(o, ", %2d", stuckKeys_memory[1]);
      $fwrite(o, ", %2d", stuckKeys_memory[2]);
      $fwrite(o, ", %2d", stuckKeys_memory[3]);
      $fwrite(o, ", %2d", stuckKeys_memory[4]);
      $fwrite(o, ", %2d", stuckKeys_memory[5]);
      $fwrite(o, ", %2d", stuckKeys_memory[6]);
      $fwrite(o, ", %2d", stuckKeys_memory[7]);
      $fwrite(o, ", %2d", stuckKeys_memory[8]);
      $fwrite(o, ", %2d", stuckKeys_memory[9]);
      $fwrite(o, ", %2d", stuckKeys_memory[10]);
      $fwrite(o, ", %2d", stuckKeys_memory[11]);
      $fwrite(o, ", %2d", stuckKeys_memory[12]);
      $fwrite(o, ", %2d", stuckKeys_memory[13]);
      $fwrite(o, ", %2d", stuckKeys_memory[14]);
      $fwrite(o, ", %2d", stuckKeys_memory[15]);
      $fwrite(o, ", %2d", stuckKeys_memory[16]);
      $fwrite(o, ", %2d", stuckKeys_memory[17]);
      $fwrite(o, ", %2d", stuckKeys_memory[18]);
      $fwrite(o, ", %2d", stuckKeys_memory[19]);
      $fwrite(o, ", %2d", stuckKeys_memory[20]);
      $fwrite(o, ", %2d", stuckKeys_memory[21]);
      $fwrite(o, ", %2d", stuckKeys_memory[22]);
      $fwrite(o, ", %2d", stuckKeys_memory[23]);
      $fwrite(o, ", %2d", stuckKeys_memory[24]);
      $fwrite(o, ", %2d", stuckKeys_memory[25]);
      $fwrite(o, ", %2d", stuckKeys_memory[26]);
      $fwrite(o, ", %2d", stuckKeys_memory[27]);
      $fwrite(o, ", %2d", stuckKeys_memory[28]);
      $fwrite(o, ", %2d", stuckKeys_memory[29]);
      $fwrite(o, ", %2d", stuckKeys_memory[30]);
      $fwrite(o, ", %2d", stuckKeys_memory[31]);
      $fwrite(o, ", %2d", stuckKeys_memory[32]);
      $fwrite(o, ", %2d", stuckKeys_memory[33]);
      $fwrite(o, ", %2d", stuckKeys_memory[34]);
      $fwrite(o, ", %2d", stuckKeys_memory[35]);
      $fwrite(o, ", %2d", stuckKeys_memory[36]);
      $fwrite(o, ", %2d", stuckKeys_memory[37]);
      $fwrite(o, ", %2d", stuckKeys_memory[38]);
      $fwrite(o, ", %2d", stuckKeys_memory[39]);
      $fwrite(o, ", %2d", stuckKeys_memory[40]);
      $fwrite(o, ", %2d", stuckKeys_memory[41]);
      $fwrite(o, ", %2d", stuckKeys_memory[42]);
      $fwrite(o, ", %2d", stuckKeys_memory[43]);
      $fwrite(o, ", %2d", stuckKeys_memory[44]);
      $fwrite(o, ", %2d", stuckKeys_memory[45]);
      $fwrite(o, ", %2d", stuckKeys_memory[46]);
      $fwrite(o, ", %2d", stuckKeys_memory[47]);
      $fwrite(o, ", %2d", stuckKeys_memory[48]);
      $fwrite(o, ", %2d", stuckKeys_memory[49]);
      $fwrite(o, ", %2d", stuckKeys_memory[50]);
      $fwrite(o, ", %2d", stuckKeys_memory[51]);
      $fwrite(o, ", %2d", stuckKeys_memory[52]);
      $fwrite(o, ", %2d", stuckKeys_memory[53]);
      $fwrite(o, ", %2d", stuckKeys_memory[54]);
      $fwrite(o, ", %2d", stuckKeys_memory[55]);
      $fwrite(o, ", %2d", stuckKeys_memory[56]);
      $fwrite(o, ", %2d", stuckKeys_memory[57]);
      $fwrite(o, ", %2d", stuckKeys_memory[58]);
      $fwrite(o, ", %2d", stuckKeys_memory[59]);
      $fwrite(o, ", %2d", stuckKeys_memory[60]);
      $fwrite(o, ", %2d", stuckKeys_memory[61]);
      $fwrite(o, ", %2d", stuckKeys_memory[62]);
      $fwrite(o, ", %2d", stuckKeys_memory[63]);
      $fwrite(o, ", %2d", stuckKeys_memory[64]);
      $fwrite(o, ", %2d", stuckKeys_memory[65]);
      $fwrite(o, ", %2d", stuckKeys_memory[66]);
      $fwrite(o, ", %2d", stuckKeys_memory[67]);
      $fwrite(o, ", %2d", stuckKeys_memory[68]);
      $fwrite(o, ", %2d", stuckKeys_memory[69]);
      $fwrite(o, ", %2d", stuckKeys_memory[70]);
      $fwrite(o, ", %2d", stuckKeys_memory[71]);
      $fwrite(o, ", %2d", stuckKeys_memory[72]);
      $fwrite(o, ", %2d", stuckKeys_memory[73]);
      $fwrite(o, ", %2d", stuckKeys_memory[74]);
      $fwrite(o, ", %2d", stuckKeys_memory[75]);
      $fwrite(o, ", %2d", stuckKeys_memory[76]);
      $fwrite(o, ", %2d", stuckKeys_memory[77]);
      $fwrite(o, ", %2d", stuckKeys_memory[78]);
      $fwrite(o, ", %2d", stuckKeys_memory[79]);
      $fwrite(o, ", %2d", stuckKeys_memory[80]);
      $fwrite(o, ", %2d", stuckKeys_memory[81]);
      $fwrite(o, ", %2d", stuckKeys_memory[82]);
      $fwrite(o, ", %2d", stuckKeys_memory[83]);
      $fwrite(o, ", %2d", stuckKeys_memory[84]);
      $fwrite(o, ", %2d", stuckKeys_memory[85]);
      $fwrite(o, ", %2d", stuckKeys_memory[86]);
      $fwrite(o, ", %2d", stuckKeys_memory[87]);
      $fwrite(o, ", %2d", stuckKeys_memory[88]);
      $fwrite(o, ", %2d", stuckKeys_memory[89]);
      $fwrite(o, ", %2d", stuckKeys_memory[90]);
      $fwrite(o, ", %2d", stuckKeys_memory[91]);
      $fwrite(o, ", %2d", stuckKeys_memory[92]);
      $fwrite(o, ", %2d", stuckKeys_memory[93]);
      $fwrite(o, ", %2d", stuckKeys_memory[94]);
      $fwrite(o, ", %2d", stuckKeys_memory[95]);
      $fwrite(o, ", %2d", stuckKeys_memory[96]);
      $fwrite(o, ", %2d", stuckKeys_memory[97]);
      $fwrite(o, ", %2d", stuckKeys_memory[98]);
      $fwrite(o, ", %2d", stuckKeys_memory[99]);
      $fwrite(o, ", %2d", stuckKeys_memory[100]);
      $fwrite(o, ", %2d", stuckKeys_memory[101]);
      $fwrite(o, ", %2d", stuckKeys_memory[102]);
      $fwrite(o, ", %2d", stuckKeys_memory[103]);
      $fwrite(o, ", %2d", stuckKeys_memory[104]);
      $fwrite(o, ", %2d", stuckKeys_memory[105]);
      $fwrite(o, ", %2d", stuckKeys_memory[106]);
      $fwrite(o, ", %2d", stuckKeys_memory[107]);
      $fwrite(o, ", %2d", stuckKeys_memory[108]);
      $fwrite(o, ", %2d", stuckKeys_memory[109]);
      $fwrite(o, ", %2d", stuckKeys_memory[110]);
      $fwrite(o, ", %2d", stuckKeys_memory[111]);
      $fwrite(o, ", %2d", stuckKeys_memory[112]);
      $fwrite(o, ", %2d", stuckKeys_memory[113]);
      $fwrite(o, ", %2d", stuckKeys_memory[114]);
      $fwrite(o, ", %2d", stuckKeys_memory[115]);
      $fwrite(o, ", %2d", stuckKeys_memory[116]);
      $fwrite(o, ", %2d", stuckKeys_memory[117]);
      $fwrite(o, ", %2d", stuckKeys_memory[118]);
      $fwrite(o, ", %2d", stuckKeys_memory[119]);
      $fwrite(o, ", %2d", stuckKeys_memory[120]);
      $fwrite(o, ", %2d", stuckKeys_memory[121]);
      $fwrite(o, ", %2d", stuckKeys_memory[122]);
      $fwrite(o, ", %2d", stuckKeys_memory[123]);
      $fwrite(o, ", %2d", stuckKeys_memory[124]);
      $fwrite(o, ", %2d", stuckKeys_memory[125]);
      $fwrite(o, ", %2d", stuckKeys_memory[126]);
      $fwrite(o, ", %2d", stuckKeys_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckKeys_1", stuckKeys_1_requestedAt, stuckKeys_1_finishedAt, stuckKeys_stuckKeys_1_returnCode, (stuckKeys_1_requestedAt > stuckKeys_1_finishedAt && stuckKeys_1_requestedAt != step), (stuckKeys_1_requestedAt < stuckKeys_1_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_1_index_20", findAndInsert_stuckKeys_1_index_20);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_0", stuckKeys_stuckKeys_1_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_1", stuckKeys_stuckKeys_1_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_2", stuckKeys_stuckKeys_1_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckKeys_stuckKeys_1_result_3", stuckKeys_stuckKeys_1_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckKeys_2", stuckKeys_2_requestedAt, stuckKeys_2_finishedAt, stuckKeys_stuckKeys_2_returnCode, (stuckKeys_2_requestedAt > stuckKeys_2_finishedAt && stuckKeys_2_requestedAt != step), (stuckKeys_2_requestedAt < stuckKeys_2_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_index_21", findAndInsert_stuckKeys_2_index_21);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_22", findAndInsert_stuckKeys_2_value_22);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_23", findAndInsert_stuckKeys_2_value_23);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_24", findAndInsert_stuckKeys_2_value_24);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckKeys_2_value_25", findAndInsert_stuckKeys_2_value_25);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 5, "stuckData", 1, stuckData_pc, stuckData_returnCode);
      $fwrite(o, "      Memory: size: %1d, width: %1d, block: %1d\n", 32, 8, 4);
      $fwrite(o, "        %2d", stuckData_memory[0]);
      $fwrite(o, ", %2d", stuckData_memory[1]);
      $fwrite(o, ", %2d", stuckData_memory[2]);
      $fwrite(o, ", %2d", stuckData_memory[3]);
      $fwrite(o, ", %2d", stuckData_memory[4]);
      $fwrite(o, ", %2d", stuckData_memory[5]);
      $fwrite(o, ", %2d", stuckData_memory[6]);
      $fwrite(o, ", %2d", stuckData_memory[7]);
      $fwrite(o, ", %2d", stuckData_memory[8]);
      $fwrite(o, ", %2d", stuckData_memory[9]);
      $fwrite(o, ", %2d", stuckData_memory[10]);
      $fwrite(o, ", %2d", stuckData_memory[11]);
      $fwrite(o, ", %2d", stuckData_memory[12]);
      $fwrite(o, ", %2d", stuckData_memory[13]);
      $fwrite(o, ", %2d", stuckData_memory[14]);
      $fwrite(o, ", %2d", stuckData_memory[15]);
      $fwrite(o, ", %2d", stuckData_memory[16]);
      $fwrite(o, ", %2d", stuckData_memory[17]);
      $fwrite(o, ", %2d", stuckData_memory[18]);
      $fwrite(o, ", %2d", stuckData_memory[19]);
      $fwrite(o, ", %2d", stuckData_memory[20]);
      $fwrite(o, ", %2d", stuckData_memory[21]);
      $fwrite(o, ", %2d", stuckData_memory[22]);
      $fwrite(o, ", %2d", stuckData_memory[23]);
      $fwrite(o, ", %2d", stuckData_memory[24]);
      $fwrite(o, ", %2d", stuckData_memory[25]);
      $fwrite(o, ", %2d", stuckData_memory[26]);
      $fwrite(o, ", %2d", stuckData_memory[27]);
      $fwrite(o, ", %2d", stuckData_memory[28]);
      $fwrite(o, ", %2d", stuckData_memory[29]);
      $fwrite(o, ", %2d", stuckData_memory[30]);
      $fwrite(o, ", %2d", stuckData_memory[31]);
      $fwrite(o, ", %2d", stuckData_memory[32]);
      $fwrite(o, ", %2d", stuckData_memory[33]);
      $fwrite(o, ", %2d", stuckData_memory[34]);
      $fwrite(o, ", %2d", stuckData_memory[35]);
      $fwrite(o, ", %2d", stuckData_memory[36]);
      $fwrite(o, ", %2d", stuckData_memory[37]);
      $fwrite(o, ", %2d", stuckData_memory[38]);
      $fwrite(o, ", %2d", stuckData_memory[39]);
      $fwrite(o, ", %2d", stuckData_memory[40]);
      $fwrite(o, ", %2d", stuckData_memory[41]);
      $fwrite(o, ", %2d", stuckData_memory[42]);
      $fwrite(o, ", %2d", stuckData_memory[43]);
      $fwrite(o, ", %2d", stuckData_memory[44]);
      $fwrite(o, ", %2d", stuckData_memory[45]);
      $fwrite(o, ", %2d", stuckData_memory[46]);
      $fwrite(o, ", %2d", stuckData_memory[47]);
      $fwrite(o, ", %2d", stuckData_memory[48]);
      $fwrite(o, ", %2d", stuckData_memory[49]);
      $fwrite(o, ", %2d", stuckData_memory[50]);
      $fwrite(o, ", %2d", stuckData_memory[51]);
      $fwrite(o, ", %2d", stuckData_memory[52]);
      $fwrite(o, ", %2d", stuckData_memory[53]);
      $fwrite(o, ", %2d", stuckData_memory[54]);
      $fwrite(o, ", %2d", stuckData_memory[55]);
      $fwrite(o, ", %2d", stuckData_memory[56]);
      $fwrite(o, ", %2d", stuckData_memory[57]);
      $fwrite(o, ", %2d", stuckData_memory[58]);
      $fwrite(o, ", %2d", stuckData_memory[59]);
      $fwrite(o, ", %2d", stuckData_memory[60]);
      $fwrite(o, ", %2d", stuckData_memory[61]);
      $fwrite(o, ", %2d", stuckData_memory[62]);
      $fwrite(o, ", %2d", stuckData_memory[63]);
      $fwrite(o, ", %2d", stuckData_memory[64]);
      $fwrite(o, ", %2d", stuckData_memory[65]);
      $fwrite(o, ", %2d", stuckData_memory[66]);
      $fwrite(o, ", %2d", stuckData_memory[67]);
      $fwrite(o, ", %2d", stuckData_memory[68]);
      $fwrite(o, ", %2d", stuckData_memory[69]);
      $fwrite(o, ", %2d", stuckData_memory[70]);
      $fwrite(o, ", %2d", stuckData_memory[71]);
      $fwrite(o, ", %2d", stuckData_memory[72]);
      $fwrite(o, ", %2d", stuckData_memory[73]);
      $fwrite(o, ", %2d", stuckData_memory[74]);
      $fwrite(o, ", %2d", stuckData_memory[75]);
      $fwrite(o, ", %2d", stuckData_memory[76]);
      $fwrite(o, ", %2d", stuckData_memory[77]);
      $fwrite(o, ", %2d", stuckData_memory[78]);
      $fwrite(o, ", %2d", stuckData_memory[79]);
      $fwrite(o, ", %2d", stuckData_memory[80]);
      $fwrite(o, ", %2d", stuckData_memory[81]);
      $fwrite(o, ", %2d", stuckData_memory[82]);
      $fwrite(o, ", %2d", stuckData_memory[83]);
      $fwrite(o, ", %2d", stuckData_memory[84]);
      $fwrite(o, ", %2d", stuckData_memory[85]);
      $fwrite(o, ", %2d", stuckData_memory[86]);
      $fwrite(o, ", %2d", stuckData_memory[87]);
      $fwrite(o, ", %2d", stuckData_memory[88]);
      $fwrite(o, ", %2d", stuckData_memory[89]);
      $fwrite(o, ", %2d", stuckData_memory[90]);
      $fwrite(o, ", %2d", stuckData_memory[91]);
      $fwrite(o, ", %2d", stuckData_memory[92]);
      $fwrite(o, ", %2d", stuckData_memory[93]);
      $fwrite(o, ", %2d", stuckData_memory[94]);
      $fwrite(o, ", %2d", stuckData_memory[95]);
      $fwrite(o, ", %2d", stuckData_memory[96]);
      $fwrite(o, ", %2d", stuckData_memory[97]);
      $fwrite(o, ", %2d", stuckData_memory[98]);
      $fwrite(o, ", %2d", stuckData_memory[99]);
      $fwrite(o, ", %2d", stuckData_memory[100]);
      $fwrite(o, ", %2d", stuckData_memory[101]);
      $fwrite(o, ", %2d", stuckData_memory[102]);
      $fwrite(o, ", %2d", stuckData_memory[103]);
      $fwrite(o, ", %2d", stuckData_memory[104]);
      $fwrite(o, ", %2d", stuckData_memory[105]);
      $fwrite(o, ", %2d", stuckData_memory[106]);
      $fwrite(o, ", %2d", stuckData_memory[107]);
      $fwrite(o, ", %2d", stuckData_memory[108]);
      $fwrite(o, ", %2d", stuckData_memory[109]);
      $fwrite(o, ", %2d", stuckData_memory[110]);
      $fwrite(o, ", %2d", stuckData_memory[111]);
      $fwrite(o, ", %2d", stuckData_memory[112]);
      $fwrite(o, ", %2d", stuckData_memory[113]);
      $fwrite(o, ", %2d", stuckData_memory[114]);
      $fwrite(o, ", %2d", stuckData_memory[115]);
      $fwrite(o, ", %2d", stuckData_memory[116]);
      $fwrite(o, ", %2d", stuckData_memory[117]);
      $fwrite(o, ", %2d", stuckData_memory[118]);
      $fwrite(o, ", %2d", stuckData_memory[119]);
      $fwrite(o, ", %2d", stuckData_memory[120]);
      $fwrite(o, ", %2d", stuckData_memory[121]);
      $fwrite(o, ", %2d", stuckData_memory[122]);
      $fwrite(o, ", %2d", stuckData_memory[123]);
      $fwrite(o, ", %2d", stuckData_memory[124]);
      $fwrite(o, ", %2d", stuckData_memory[125]);
      $fwrite(o, ", %2d", stuckData_memory[126]);
      $fwrite(o, ", %2d", stuckData_memory[127]);
      $fwrite(o, "\n");
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);
      $fwrite(o, "      Transactions:\n");
      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "get", "stuckData_3", stuckData_3_requestedAt, stuckData_3_finishedAt, stuckData_stuckData_3_returnCode, (stuckData_3_requestedAt > stuckData_3_finishedAt && stuckData_3_requestedAt != step), (stuckData_3_requestedAt < stuckData_3_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_3_index_26", findAndInsert_stuckData_3_index_26);

      $fwrite(o, "          Outputs     :\n");

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_0", stuckData_stuckData_3_result_0);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_1", stuckData_stuckData_3_result_1);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_2", stuckData_stuckData_3_result_2);

      $fwrite(o, "            %-38s = %1d\n", "stuckData_stuckData_3_result_3", stuckData_stuckData_3_result_3);

      $fwrite(o, "        Transaction   : %-8s - %-16s  requested at: %1d, finished at: %1d, returnCode: %1d, executable: %1d, finished: %1d\n", "set", "stuckData_4", stuckData_4_requestedAt, stuckData_4_finishedAt, stuckData_stuckData_4_returnCode, (stuckData_4_requestedAt > stuckData_4_finishedAt && stuckData_4_requestedAt != step), (stuckData_4_requestedAt < stuckData_4_finishedAt));

      $fwrite(o, "          Inputs      :\n");
      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_index_27", findAndInsert_stuckData_4_index_27);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_28", findAndInsert_stuckData_4_value_28);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_29", findAndInsert_stuckData_4_value_29);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_30", findAndInsert_stuckData_4_value_30);

      $fwrite(o, "            %-38s = %1d\n", "findAndInsert_stuckData_4_value_31", findAndInsert_stuckData_4_value_31);

      $fwrite(o, "    Process: %1d - %-21s instructions: %1d, pc: %1d, rc: %1d\n", 6, "findAndInsert", 53, findAndInsert_pc, findAndInsert_returnCode);
      $fwrite(o, "      Registers :\n");
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_0", findAndInsert_index_0);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_1", findAndInsert_size_1);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_2", findAndInsert_isLeaf_2);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_3", findAndInsert_nextFree_3);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_4", findAndInsert_Key_0_4);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_5", findAndInsert_KeyCompares_0_5);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_6", findAndInsert_KeyCollapse_0_6);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_7", findAndInsert_Data_0_7);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_8", findAndInsert_Key_1_8);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_9", findAndInsert_KeyCompares_1_9);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_10", findAndInsert_KeyCollapse_1_10);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_11", findAndInsert_Data_1_11);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_12", findAndInsert_Key_2_12);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_13", findAndInsert_KeyCompares_2_13);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_14", findAndInsert_KeyCollapse_2_14);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_15", findAndInsert_Data_2_15);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_16", findAndInsert_Key_3_16);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_17", findAndInsert_KeyCompares_3_17);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_18", findAndInsert_KeyCollapse_3_18);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_19", findAndInsert_Data_3_19);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_1_index_20", findAndInsert_stuckKeys_1_index_20);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_index_21", findAndInsert_stuckKeys_2_index_21);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_22", findAndInsert_stuckKeys_2_value_22);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_23", findAndInsert_stuckKeys_2_value_23);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_24", findAndInsert_stuckKeys_2_value_24);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckKeys_2_value_25", findAndInsert_stuckKeys_2_value_25);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_3_index_26", findAndInsert_stuckData_3_index_26);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_index_27", findAndInsert_stuckData_4_index_27);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_28", findAndInsert_stuckData_4_value_28);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_29", findAndInsert_stuckData_4_value_29);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_30", findAndInsert_stuckData_4_value_30);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckData_4_value_31", findAndInsert_stuckData_4_value_31);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckSize_5_index_32", findAndInsert_stuckSize_5_index_32);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckSize_6_index_33", findAndInsert_stuckSize_6_index_33);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckSize_6_value_34", findAndInsert_stuckSize_6_value_34);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsLeaf_7_index_35", findAndInsert_stuckIsLeaf_7_index_35);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsLeaf_8_index_36", findAndInsert_stuckIsLeaf_8_index_36);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsLeaf_8_value_37", findAndInsert_stuckIsLeaf_8_value_37);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_38", findAndInsert_Found_38);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_39", findAndInsert_Key_39);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_40", findAndInsert_FoundKey_40);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_41", findAndInsert_Data_41);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_42", findAndInsert_BtreeIndex_42);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_43", findAndInsert_StuckIndex_43);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_44", findAndInsert_MergeSuccess_44);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_i_45", findAndInsert_i_45);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_j_46", findAndInsert_j_46);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_47", findAndInsert_index_47);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_48", findAndInsert_size_48);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_49", findAndInsert_isLeaf_49);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_50", findAndInsert_nextFree_50);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_51", findAndInsert_Key_0_51);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_52", findAndInsert_KeyCompares_0_52);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_53", findAndInsert_KeyCollapse_0_53);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_54", findAndInsert_Data_0_54);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_55", findAndInsert_Key_1_55);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_56", findAndInsert_KeyCompares_1_56);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_57", findAndInsert_KeyCollapse_1_57);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_58", findAndInsert_Data_1_58);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_59", findAndInsert_Key_2_59);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_60", findAndInsert_KeyCompares_2_60);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_61", findAndInsert_KeyCollapse_2_61);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_62", findAndInsert_Data_2_62);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_63", findAndInsert_Key_3_63);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_64", findAndInsert_KeyCompares_3_64);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_65", findAndInsert_KeyCollapse_3_65);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_66", findAndInsert_Data_3_66);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_67", findAndInsert_Found_67);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_68", findAndInsert_Key_68);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_69", findAndInsert_FoundKey_69);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_70", findAndInsert_Data_70);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_71", findAndInsert_BtreeIndex_71);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_72", findAndInsert_StuckIndex_72);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_73", findAndInsert_MergeSuccess_73);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_74", findAndInsert_index_74);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_75", findAndInsert_size_75);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_76", findAndInsert_isLeaf_76);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_77", findAndInsert_nextFree_77);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_78", findAndInsert_Key_0_78);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_79", findAndInsert_KeyCompares_0_79);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_80", findAndInsert_KeyCollapse_0_80);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_81", findAndInsert_Data_0_81);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_82", findAndInsert_Key_1_82);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_83", findAndInsert_KeyCompares_1_83);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_84", findAndInsert_KeyCollapse_1_84);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_85", findAndInsert_Data_1_85);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_86", findAndInsert_Key_2_86);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_87", findAndInsert_KeyCompares_2_87);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_88", findAndInsert_KeyCollapse_2_88);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_89", findAndInsert_Data_2_89);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_90", findAndInsert_Key_3_90);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_91", findAndInsert_KeyCompares_3_91);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_92", findAndInsert_KeyCollapse_3_92);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_93", findAndInsert_Data_3_93);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_94", findAndInsert_Found_94);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_95", findAndInsert_Key_95);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_96", findAndInsert_FoundKey_96);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_97", findAndInsert_Data_97);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_98", findAndInsert_BtreeIndex_98);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_99", findAndInsert_StuckIndex_99);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_100", findAndInsert_MergeSuccess_100);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_101", findAndInsert_index_101);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_102", findAndInsert_size_102);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_103", findAndInsert_isLeaf_103);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_104", findAndInsert_nextFree_104);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_105", findAndInsert_Key_0_105);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_106", findAndInsert_KeyCompares_0_106);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_107", findAndInsert_KeyCollapse_0_107);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_108", findAndInsert_Data_0_108);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_109", findAndInsert_Key_1_109);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_110", findAndInsert_KeyCompares_1_110);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_111", findAndInsert_KeyCollapse_1_111);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_112", findAndInsert_Data_1_112);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_113", findAndInsert_Key_2_113);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_114", findAndInsert_KeyCompares_2_114);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_115", findAndInsert_KeyCollapse_2_115);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_116", findAndInsert_Data_2_116);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_117", findAndInsert_Key_3_117);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_118", findAndInsert_KeyCompares_3_118);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_119", findAndInsert_KeyCollapse_3_119);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_120", findAndInsert_Data_3_120);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_121", findAndInsert_Found_121);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_122", findAndInsert_Key_122);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_123", findAndInsert_FoundKey_123);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_124", findAndInsert_Data_124);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_125", findAndInsert_BtreeIndex_125);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_126", findAndInsert_StuckIndex_126);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_127", findAndInsert_MergeSuccess_127);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_128", findAndInsert_index_128);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_129", findAndInsert_size_129);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_130", findAndInsert_isLeaf_130);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_131", findAndInsert_nextFree_131);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_132", findAndInsert_Key_0_132);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_133", findAndInsert_KeyCompares_0_133);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_134", findAndInsert_KeyCollapse_0_134);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_135", findAndInsert_Data_0_135);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_136", findAndInsert_Key_1_136);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_137", findAndInsert_KeyCompares_1_137);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_138", findAndInsert_KeyCollapse_1_138);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_139", findAndInsert_Data_1_139);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_140", findAndInsert_Key_2_140);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_141", findAndInsert_KeyCompares_2_141);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_142", findAndInsert_KeyCollapse_2_142);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_143", findAndInsert_Data_2_143);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_144", findAndInsert_Key_3_144);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_145", findAndInsert_KeyCompares_3_145);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_146", findAndInsert_KeyCollapse_3_146);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_147", findAndInsert_Data_3_147);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_148", findAndInsert_Found_148);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_149", findAndInsert_Key_149);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_150", findAndInsert_FoundKey_150);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_151", findAndInsert_Data_151);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_152", findAndInsert_BtreeIndex_152);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_153", findAndInsert_StuckIndex_153);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_154", findAndInsert_MergeSuccess_154);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childKey_155", findAndInsert_childKey_155);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childData_156", findAndInsert_childData_156);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexLeft_157", findAndInsert_indexLeft_157);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexRight_158", findAndInsert_indexRight_158);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_midKey_159", findAndInsert_midKey_159);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_freeNext_9_index_160", findAndInsert_freeNext_9_index_160);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_freeNext_10_index_161", findAndInsert_freeNext_10_index_161);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_freeNext_10_value_162", findAndInsert_freeNext_10_value_162);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsFree_11_index_163", findAndInsert_stuckIsFree_11_index_163);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_stuckIsFree_11_value_164", findAndInsert_stuckIsFree_11_value_164);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_root_165", findAndInsert_root_165);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_next_166", findAndInsert_next_166);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_167", findAndInsert_isLeaf_167);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isFree_168", findAndInsert_isFree_168);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_169", findAndInsert_index_169);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_170", findAndInsert_size_170);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_171", findAndInsert_isLeaf_171);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_172", findAndInsert_nextFree_172);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_173", findAndInsert_Key_0_173);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_174", findAndInsert_KeyCompares_0_174);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_175", findAndInsert_KeyCollapse_0_175);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_176", findAndInsert_Data_0_176);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_177", findAndInsert_Key_1_177);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_178", findAndInsert_KeyCompares_1_178);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_179", findAndInsert_KeyCollapse_1_179);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_180", findAndInsert_Data_1_180);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_181", findAndInsert_Key_2_181);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_182", findAndInsert_KeyCompares_2_182);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_183", findAndInsert_KeyCollapse_2_183);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_184", findAndInsert_Data_2_184);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_185", findAndInsert_Key_3_185);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_186", findAndInsert_KeyCompares_3_186);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_187", findAndInsert_KeyCollapse_3_187);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_188", findAndInsert_Data_3_188);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_189", findAndInsert_Found_189);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_190", findAndInsert_Key_190);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_191", findAndInsert_FoundKey_191);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_192", findAndInsert_Data_192);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_193", findAndInsert_BtreeIndex_193);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_194", findAndInsert_StuckIndex_194);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_195", findAndInsert_MergeSuccess_195);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_index_196", findAndInsert_index_196);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_197", findAndInsert_size_197);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isLeaf_198", findAndInsert_isLeaf_198);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_nextFree_199", findAndInsert_nextFree_199);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_0_200", findAndInsert_Key_0_200);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_0_201", findAndInsert_KeyCompares_0_201);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_0_202", findAndInsert_KeyCollapse_0_202);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_0_203", findAndInsert_Data_0_203);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_1_204", findAndInsert_Key_1_204);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_1_205", findAndInsert_KeyCompares_1_205);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_1_206", findAndInsert_KeyCollapse_1_206);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_1_207", findAndInsert_Data_1_207);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_2_208", findAndInsert_Key_2_208);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_2_209", findAndInsert_KeyCompares_2_209);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_2_210", findAndInsert_KeyCollapse_2_210);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_2_211", findAndInsert_Data_2_211);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_3_212", findAndInsert_Key_3_212);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCompares_3_213", findAndInsert_KeyCompares_3_213);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_KeyCollapse_3_214", findAndInsert_KeyCollapse_3_214);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_3_215", findAndInsert_Data_3_215);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Found_216", findAndInsert_Found_216);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Key_217", findAndInsert_Key_217);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_FoundKey_218", findAndInsert_FoundKey_218);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_Data_219", findAndInsert_Data_219);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_BtreeIndex_220", findAndInsert_BtreeIndex_220);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_StuckIndex_221", findAndInsert_StuckIndex_221);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_MergeSuccess_222", findAndInsert_MergeSuccess_222);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childKey_223", findAndInsert_childKey_223);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_size_224", findAndInsert_size_224);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_childData_225", findAndInsert_childData_225);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexLeft_226", findAndInsert_indexLeft_226);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_indexRight_227", findAndInsert_indexRight_227);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_midKey_228", findAndInsert_midKey_228);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_success_229", findAndInsert_success_229);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_test_230", findAndInsert_test_230);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_next_231", findAndInsert_next_231);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_root_232", findAndInsert_root_232);
      $fwrite(o, "        Register: %-32s = %1d\n",  "findAndInsert_isFree_233", findAndInsert_isFree_233);
      $fclose(o);
    end
  endtask
endmodule
